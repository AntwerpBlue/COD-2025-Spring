
`timescale 1ns/1ps
module mem_bram #(
    parameter ADDR_WIDTH = 10,		//地址宽度
    parameter DATA_WIDTH = 128		//数据宽度
)(
    input                   clk,   // Clock
    input [ADDR_WIDTH-1:0]  raddr,  // Address
    input [ADDR_WIDTH-1:0]  waddr,  // Address
    input [DATA_WIDTH-1:0]  din,   // Data Input
    input                   we,    // Write Enable
    output [DATA_WIDTH-1:0] dout   // Data Output
); 
    reg [ADDR_WIDTH-1:0] addr_r;  // Address Register
    reg [DATA_WIDTH-1:0] ram [0:(1 << ADDR_WIDTH)-1];
    integer i;
    initial begin
        ram[0][31:0] = 32'd1870585436;
        ram[0][63:32] = 32'd2069472944;
        ram[0][95:64] = 32'd861516427;
        ram[0][127:96] = 32'd3350406635;
        ram[1][31:0] = 32'd1555224870;
        ram[1][63:32] = 32'd2154190107;
        ram[1][95:64] = 32'd1402063009;
        ram[1][127:96] = 32'd2041861951;
        ram[2][31:0] = 32'd3505230681;
        ram[2][63:32] = 32'd1323063753;
        ram[2][95:64] = 32'd4271687727;
        ram[2][127:96] = 32'd2298463057;
        ram[3][31:0] = 32'd1768449257;
        ram[3][63:32] = 32'd4162140124;
        ram[3][95:64] = 32'd539032534;
        ram[3][127:96] = 32'd1119003857;
        ram[4][31:0] = 32'd3925987810;
        ram[4][63:32] = 32'd1949417226;
        ram[4][95:64] = 32'd1569000094;
        ram[4][127:96] = 32'd1070811302;
        ram[5][31:0] = 32'd592586045;
        ram[5][63:32] = 32'd10047926;
        ram[5][95:64] = 32'd1621961986;
        ram[5][127:96] = 32'd2945448156;
        ram[6][31:0] = 32'd2159349817;
        ram[6][63:32] = 32'd1147999157;
        ram[6][95:64] = 32'd1486386312;
        ram[6][127:96] = 32'd1798709310;
        ram[7][31:0] = 32'd4030679079;
        ram[7][63:32] = 32'd3629881189;
        ram[7][95:64] = 32'd1193996624;
        ram[7][127:96] = 32'd3527005491;
        ram[8][31:0] = 32'd3844512050;
        ram[8][63:32] = 32'd1146315537;
        ram[8][95:64] = 32'd1289644746;
        ram[8][127:96] = 32'd1604560142;
        ram[9][31:0] = 32'd1757996162;
        ram[9][63:32] = 32'd3077452828;
        ram[9][95:64] = 32'd179744430;
        ram[9][127:96] = 32'd2872399735;
        ram[10][31:0] = 32'd1444412845;
        ram[10][63:32] = 32'd660859156;
        ram[10][95:64] = 32'd3414355641;
        ram[10][127:96] = 32'd3210668433;
        ram[11][31:0] = 32'd1380847095;
        ram[11][63:32] = 32'd2933273070;
        ram[11][95:64] = 32'd1882782061;
        ram[11][127:96] = 32'd999277383;
        ram[12][31:0] = 32'd2577690104;
        ram[12][63:32] = 32'd2828154457;
        ram[12][95:64] = 32'd3713624851;
        ram[12][127:96] = 32'd3352351002;
        ram[13][31:0] = 32'd3291818831;
        ram[13][63:32] = 32'd48823010;
        ram[13][95:64] = 32'd1614540136;
        ram[13][127:96] = 32'd4041042842;
        ram[14][31:0] = 32'd2473651066;
        ram[14][63:32] = 32'd400692079;
        ram[14][95:64] = 32'd2831688436;
        ram[14][127:96] = 32'd1487397129;
        ram[15][31:0] = 32'd3735645991;
        ram[15][63:32] = 32'd3519769342;
        ram[15][95:64] = 32'd504570280;
        ram[15][127:96] = 32'd2384061833;
        ram[16][31:0] = 32'd4168218661;
        ram[16][63:32] = 32'd3399266989;
        ram[16][95:64] = 32'd876819121;
        ram[16][127:96] = 32'd2886172558;
        ram[17][31:0] = 32'd3542550272;
        ram[17][63:32] = 32'd3387089861;
        ram[17][95:64] = 32'd3874690545;
        ram[17][127:96] = 32'd963159638;
        ram[18][31:0] = 32'd3699586661;
        ram[18][63:32] = 32'd297754104;
        ram[18][95:64] = 32'd3146623705;
        ram[18][127:96] = 32'd3972422453;
        ram[19][31:0] = 32'd1051232611;
        ram[19][63:32] = 32'd998193764;
        ram[19][95:64] = 32'd3095344887;
        ram[19][127:96] = 32'd466432104;
        ram[20][31:0] = 32'd3440150321;
        ram[20][63:32] = 32'd2716768050;
        ram[20][95:64] = 32'd979668869;
        ram[20][127:96] = 32'd2260163579;
        ram[21][31:0] = 32'd1958613062;
        ram[21][63:32] = 32'd3703089126;
        ram[21][95:64] = 32'd623629618;
        ram[21][127:96] = 32'd3303907992;
        ram[22][31:0] = 32'd1506464650;
        ram[22][63:32] = 32'd1036241526;
        ram[22][95:64] = 32'd548807498;
        ram[22][127:96] = 32'd3415150818;
        ram[23][31:0] = 32'd4105109197;
        ram[23][63:32] = 32'd4048368480;
        ram[23][95:64] = 32'd2640578934;
        ram[23][127:96] = 32'd411761706;
        ram[24][31:0] = 32'd1607774016;
        ram[24][63:32] = 32'd2681259618;
        ram[24][95:64] = 32'd1885671812;
        ram[24][127:96] = 32'd2668054470;
        ram[25][31:0] = 32'd3329548407;
        ram[25][63:32] = 32'd293268391;
        ram[25][95:64] = 32'd3476251709;
        ram[25][127:96] = 32'd3105134583;
        ram[26][31:0] = 32'd1835365570;
        ram[26][63:32] = 32'd1914703890;
        ram[26][95:64] = 32'd3973347769;
        ram[26][127:96] = 32'd2329785644;
        ram[27][31:0] = 32'd61872566;
        ram[27][63:32] = 32'd2828290416;
        ram[27][95:64] = 32'd1786256609;
        ram[27][127:96] = 32'd2224133112;
        ram[28][31:0] = 32'd2138465740;
        ram[28][63:32] = 32'd2509755899;
        ram[28][95:64] = 32'd759874881;
        ram[28][127:96] = 32'd1862517686;
        ram[29][31:0] = 32'd1148833960;
        ram[29][63:32] = 32'd1057530362;
        ram[29][95:64] = 32'd2857138427;
        ram[29][127:96] = 32'd2989373656;
        ram[30][31:0] = 32'd132670189;
        ram[30][63:32] = 32'd371426538;
        ram[30][95:64] = 32'd1367201542;
        ram[30][127:96] = 32'd2458710516;
        ram[31][31:0] = 32'd1496960271;
        ram[31][63:32] = 32'd1825838587;
        ram[31][95:64] = 32'd3622232671;
        ram[31][127:96] = 32'd415964961;
        ram[32][31:0] = 32'd3976736584;
        ram[32][63:32] = 32'd1885285401;
        ram[32][95:64] = 32'd454112648;
        ram[32][127:96] = 32'd351680695;
        ram[33][31:0] = 32'd4027336748;
        ram[33][63:32] = 32'd1549772363;
        ram[33][95:64] = 32'd167479484;
        ram[33][127:96] = 32'd1960021159;
        ram[34][31:0] = 32'd3552771192;
        ram[34][63:32] = 32'd3115074711;
        ram[34][95:64] = 32'd2291202182;
        ram[34][127:96] = 32'd598541164;
        ram[35][31:0] = 32'd684175502;
        ram[35][63:32] = 32'd3385276041;
        ram[35][95:64] = 32'd720488543;
        ram[35][127:96] = 32'd1761678698;
        ram[36][31:0] = 32'd725755827;
        ram[36][63:32] = 32'd2276121759;
        ram[36][95:64] = 32'd1978812597;
        ram[36][127:96] = 32'd3498313420;
        ram[37][31:0] = 32'd2210961168;
        ram[37][63:32] = 32'd404226320;
        ram[37][95:64] = 32'd1729930243;
        ram[37][127:96] = 32'd302678610;
        ram[38][31:0] = 32'd422264761;
        ram[38][63:32] = 32'd352254805;
        ram[38][95:64] = 32'd1437003575;
        ram[38][127:96] = 32'd979919250;
        ram[39][31:0] = 32'd1698941605;
        ram[39][63:32] = 32'd1981510702;
        ram[39][95:64] = 32'd2395849516;
        ram[39][127:96] = 32'd4008254182;
        ram[40][31:0] = 32'd2220794859;
        ram[40][63:32] = 32'd2656187847;
        ram[40][95:64] = 32'd775522268;
        ram[40][127:96] = 32'd3495425455;
        ram[41][31:0] = 32'd2460820341;
        ram[41][63:32] = 32'd3760476342;
        ram[41][95:64] = 32'd1889795081;
        ram[41][127:96] = 32'd3268472177;
        ram[42][31:0] = 32'd2286702594;
        ram[42][63:32] = 32'd1140743891;
        ram[42][95:64] = 32'd3539743854;
        ram[42][127:96] = 32'd3511614128;
        ram[43][31:0] = 32'd2616985559;
        ram[43][63:32] = 32'd422894365;
        ram[43][95:64] = 32'd3085808268;
        ram[43][127:96] = 32'd3567745488;
        ram[44][31:0] = 32'd643849309;
        ram[44][63:32] = 32'd2295881178;
        ram[44][95:64] = 32'd2677761729;
        ram[44][127:96] = 32'd2886227464;
        ram[45][31:0] = 32'd1980496809;
        ram[45][63:32] = 32'd3424920418;
        ram[45][95:64] = 32'd1222529405;
        ram[45][127:96] = 32'd4192569996;
        ram[46][31:0] = 32'd961772350;
        ram[46][63:32] = 32'd767163713;
        ram[46][95:64] = 32'd862037870;
        ram[46][127:96] = 32'd3131077888;
        ram[47][31:0] = 32'd1685919072;
        ram[47][63:32] = 32'd133639369;
        ram[47][95:64] = 32'd4284820396;
        ram[47][127:96] = 32'd1124573723;
        ram[48][31:0] = 32'd597630141;
        ram[48][63:32] = 32'd2053860581;
        ram[48][95:64] = 32'd2242595831;
        ram[48][127:96] = 32'd186646160;
        ram[49][31:0] = 32'd2562666729;
        ram[49][63:32] = 32'd4294944672;
        ram[49][95:64] = 32'd1771443269;
        ram[49][127:96] = 32'd1445264864;
        ram[50][31:0] = 32'd3635105000;
        ram[50][63:32] = 32'd2051129310;
        ram[50][95:64] = 32'd4173384693;
        ram[50][127:96] = 32'd1663091370;
        ram[51][31:0] = 32'd3125904639;
        ram[51][63:32] = 32'd349509858;
        ram[51][95:64] = 32'd871555750;
        ram[51][127:96] = 32'd3823761644;
        ram[52][31:0] = 32'd3010632164;
        ram[52][63:32] = 32'd885491266;
        ram[52][95:64] = 32'd2556735740;
        ram[52][127:96] = 32'd3337632621;
        ram[53][31:0] = 32'd4150766495;
        ram[53][63:32] = 32'd371999850;
        ram[53][95:64] = 32'd3364977113;
        ram[53][127:96] = 32'd2179149214;
        ram[54][31:0] = 32'd2231833515;
        ram[54][63:32] = 32'd797224449;
        ram[54][95:64] = 32'd2791150383;
        ram[54][127:96] = 32'd393784553;
        ram[55][31:0] = 32'd4233481341;
        ram[55][63:32] = 32'd285286831;
        ram[55][95:64] = 32'd4222144713;
        ram[55][127:96] = 32'd308136402;
        ram[56][31:0] = 32'd3721336189;
        ram[56][63:32] = 32'd4158612666;
        ram[56][95:64] = 32'd326705489;
        ram[56][127:96] = 32'd4147188654;
        ram[57][31:0] = 32'd3918629529;
        ram[57][63:32] = 32'd3264330583;
        ram[57][95:64] = 32'd1100096081;
        ram[57][127:96] = 32'd1221449456;
        ram[58][31:0] = 32'd4110523392;
        ram[58][63:32] = 32'd2577766004;
        ram[58][95:64] = 32'd1597413610;
        ram[58][127:96] = 32'd1995153683;
        ram[59][31:0] = 32'd3308823479;
        ram[59][63:32] = 32'd3710833553;
        ram[59][95:64] = 32'd1412625860;
        ram[59][127:96] = 32'd808220211;
        ram[60][31:0] = 32'd2785262700;
        ram[60][63:32] = 32'd3647911902;
        ram[60][95:64] = 32'd1066521417;
        ram[60][127:96] = 32'd488961057;
        ram[61][31:0] = 32'd2896346636;
        ram[61][63:32] = 32'd2801824671;
        ram[61][95:64] = 32'd2321687399;
        ram[61][127:96] = 32'd2088915050;
        ram[62][31:0] = 32'd2567675747;
        ram[62][63:32] = 32'd634363534;
        ram[62][95:64] = 32'd3563604010;
        ram[62][127:96] = 32'd528276894;
        ram[63][31:0] = 32'd3233104755;
        ram[63][63:32] = 32'd2251486923;
        ram[63][95:64] = 32'd4129721780;
        ram[63][127:96] = 32'd4293329829;
        ram[64][31:0] = 32'd214161842;
        ram[64][63:32] = 32'd2962833118;
        ram[64][95:64] = 32'd3768261454;
        ram[64][127:96] = 32'd735052196;
        ram[65][31:0] = 32'd2209658087;
        ram[65][63:32] = 32'd2908678289;
        ram[65][95:64] = 32'd3668048787;
        ram[65][127:96] = 32'd2095898228;
        ram[66][31:0] = 32'd1563802891;
        ram[66][63:32] = 32'd2676695456;
        ram[66][95:64] = 32'd247106196;
        ram[66][127:96] = 32'd1193893598;
        ram[67][31:0] = 32'd458908171;
        ram[67][63:32] = 32'd3243925981;
        ram[67][95:64] = 32'd1805982290;
        ram[67][127:96] = 32'd2912190139;
        ram[68][31:0] = 32'd495494873;
        ram[68][63:32] = 32'd793232809;
        ram[68][95:64] = 32'd1240901263;
        ram[68][127:96] = 32'd94646178;
        ram[69][31:0] = 32'd3369498205;
        ram[69][63:32] = 32'd76492403;
        ram[69][95:64] = 32'd3087657609;
        ram[69][127:96] = 32'd1301179723;
        ram[70][31:0] = 32'd535207050;
        ram[70][63:32] = 32'd866061806;
        ram[70][95:64] = 32'd1396158732;
        ram[70][127:96] = 32'd4134955926;
        ram[71][31:0] = 32'd1470833253;
        ram[71][63:32] = 32'd531515270;
        ram[71][95:64] = 32'd1109364526;
        ram[71][127:96] = 32'd2077233220;
        ram[72][31:0] = 32'd3761039539;
        ram[72][63:32] = 32'd940573815;
        ram[72][95:64] = 32'd1919999915;
        ram[72][127:96] = 32'd2648754452;
        ram[73][31:0] = 32'd3646512956;
        ram[73][63:32] = 32'd120765790;
        ram[73][95:64] = 32'd2294789991;
        ram[73][127:96] = 32'd431105951;
        ram[74][31:0] = 32'd1128855117;
        ram[74][63:32] = 32'd4171669338;
        ram[74][95:64] = 32'd3316398040;
        ram[74][127:96] = 32'd1285349339;
        ram[75][31:0] = 32'd4260493041;
        ram[75][63:32] = 32'd779647779;
        ram[75][95:64] = 32'd2759854552;
        ram[75][127:96] = 32'd3371624447;
        ram[76][31:0] = 32'd2015865801;
        ram[76][63:32] = 32'd1517077955;
        ram[76][95:64] = 32'd1400119106;
        ram[76][127:96] = 32'd3130498011;
        ram[77][31:0] = 32'd2611705428;
        ram[77][63:32] = 32'd3941608837;
        ram[77][95:64] = 32'd3094631771;
        ram[77][127:96] = 32'd1449524691;
        ram[78][31:0] = 32'd240548675;
        ram[78][63:32] = 32'd402285906;
        ram[78][95:64] = 32'd3194236288;
        ram[78][127:96] = 32'd3309303920;
        ram[79][31:0] = 32'd838957123;
        ram[79][63:32] = 32'd3819728146;
        ram[79][95:64] = 32'd530093518;
        ram[79][127:96] = 32'd700414460;
        ram[80][31:0] = 32'd1447166892;
        ram[80][63:32] = 32'd4078285937;
        ram[80][95:64] = 32'd4172724571;
        ram[80][127:96] = 32'd2407757486;
        ram[81][31:0] = 32'd1292645181;
        ram[81][63:32] = 32'd2757063505;
        ram[81][95:64] = 32'd3024984000;
        ram[81][127:96] = 32'd318989378;
        ram[82][31:0] = 32'd3131202390;
        ram[82][63:32] = 32'd2281836126;
        ram[82][95:64] = 32'd1703867803;
        ram[82][127:96] = 32'd2887064224;
        ram[83][31:0] = 32'd3238606923;
        ram[83][63:32] = 32'd4014888690;
        ram[83][95:64] = 32'd1647084470;
        ram[83][127:96] = 32'd115410482;
        ram[84][31:0] = 32'd2188727585;
        ram[84][63:32] = 32'd325795203;
        ram[84][95:64] = 32'd3556465203;
        ram[84][127:96] = 32'd2720908177;
        ram[85][31:0] = 32'd1208493341;
        ram[85][63:32] = 32'd829190514;
        ram[85][95:64] = 32'd2723057950;
        ram[85][127:96] = 32'd1424482524;
        ram[86][31:0] = 32'd281373290;
        ram[86][63:32] = 32'd3249490296;
        ram[86][95:64] = 32'd3397465739;
        ram[86][127:96] = 32'd184952467;
        ram[87][31:0] = 32'd3476652391;
        ram[87][63:32] = 32'd2061620473;
        ram[87][95:64] = 32'd2859227479;
        ram[87][127:96] = 32'd844257886;
        ram[88][31:0] = 32'd147931898;
        ram[88][63:32] = 32'd1647595599;
        ram[88][95:64] = 32'd3966319412;
        ram[88][127:96] = 32'd529744175;
        ram[89][31:0] = 32'd3033278383;
        ram[89][63:32] = 32'd1970531824;
        ram[89][95:64] = 32'd928067253;
        ram[89][127:96] = 32'd4082684122;
        ram[90][31:0] = 32'd1883443685;
        ram[90][63:32] = 32'd1749764396;
        ram[90][95:64] = 32'd3612932426;
        ram[90][127:96] = 32'd3770020475;
        ram[91][31:0] = 32'd4047546126;
        ram[91][63:32] = 32'd2422224454;
        ram[91][95:64] = 32'd2115114658;
        ram[91][127:96] = 32'd695560474;
        ram[92][31:0] = 32'd3673022184;
        ram[92][63:32] = 32'd3255881668;
        ram[92][95:64] = 32'd1599783578;
        ram[92][127:96] = 32'd1555706204;
        ram[93][31:0] = 32'd3348876813;
        ram[93][63:32] = 32'd6943526;
        ram[93][95:64] = 32'd1975409823;
        ram[93][127:96] = 32'd137070870;
        ram[94][31:0] = 32'd3383574487;
        ram[94][63:32] = 32'd258678087;
        ram[94][95:64] = 32'd1707274193;
        ram[94][127:96] = 32'd76696075;
        ram[95][31:0] = 32'd4157069748;
        ram[95][63:32] = 32'd3760007301;
        ram[95][95:64] = 32'd1718641206;
        ram[95][127:96] = 32'd2799539366;
        ram[96][31:0] = 32'd2543455748;
        ram[96][63:32] = 32'd2580136147;
        ram[96][95:64] = 32'd2578070289;
        ram[96][127:96] = 32'd2510655191;
        ram[97][31:0] = 32'd2217298716;
        ram[97][63:32] = 32'd2233888802;
        ram[97][95:64] = 32'd1776181937;
        ram[97][127:96] = 32'd4156755592;
        ram[98][31:0] = 32'd4188547242;
        ram[98][63:32] = 32'd584673643;
        ram[98][95:64] = 32'd1695524531;
        ram[98][127:96] = 32'd1000866044;
        ram[99][31:0] = 32'd179786261;
        ram[99][63:32] = 32'd1048663066;
        ram[99][95:64] = 32'd498624505;
        ram[99][127:96] = 32'd3647612275;
        ram[100][31:0] = 32'd3091846241;
        ram[100][63:32] = 32'd1021537005;
        ram[100][95:64] = 32'd246986956;
        ram[100][127:96] = 32'd1922485250;
        ram[101][31:0] = 32'd284306586;
        ram[101][63:32] = 32'd411101395;
        ram[101][95:64] = 32'd2569288348;
        ram[101][127:96] = 32'd1877487673;
        ram[102][31:0] = 32'd543094332;
        ram[102][63:32] = 32'd2882373882;
        ram[102][95:64] = 32'd3422075366;
        ram[102][127:96] = 32'd2049410600;
        ram[103][31:0] = 32'd35661170;
        ram[103][63:32] = 32'd2121687939;
        ram[103][95:64] = 32'd3438809741;
        ram[103][127:96] = 32'd2824809495;
        ram[104][31:0] = 32'd3861098664;
        ram[104][63:32] = 32'd3832011826;
        ram[104][95:64] = 32'd1591263160;
        ram[104][127:96] = 32'd188335908;
        ram[105][31:0] = 32'd3279180000;
        ram[105][63:32] = 32'd3567358548;
        ram[105][95:64] = 32'd2973342047;
        ram[105][127:96] = 32'd3889544275;
        ram[106][31:0] = 32'd458707520;
        ram[106][63:32] = 32'd1849732206;
        ram[106][95:64] = 32'd138557177;
        ram[106][127:96] = 32'd1979928705;
        ram[107][31:0] = 32'd1479974522;
        ram[107][63:32] = 32'd3385333427;
        ram[107][95:64] = 32'd2489047385;
        ram[107][127:96] = 32'd723449661;
        ram[108][31:0] = 32'd1474827311;
        ram[108][63:32] = 32'd1227238690;
        ram[108][95:64] = 32'd3881600915;
        ram[108][127:96] = 32'd1781223650;
        ram[109][31:0] = 32'd1024435444;
        ram[109][63:32] = 32'd2319963295;
        ram[109][95:64] = 32'd3957892093;
        ram[109][127:96] = 32'd1018885802;
        ram[110][31:0] = 32'd118271122;
        ram[110][63:32] = 32'd3910731565;
        ram[110][95:64] = 32'd3875418356;
        ram[110][127:96] = 32'd2309805798;
        ram[111][31:0] = 32'd3460837510;
        ram[111][63:32] = 32'd57979874;
        ram[111][95:64] = 32'd185249361;
        ram[111][127:96] = 32'd560305466;
        ram[112][31:0] = 32'd4199406484;
        ram[112][63:32] = 32'd2000661367;
        ram[112][95:64] = 32'd1220832376;
        ram[112][127:96] = 32'd2278524113;
        ram[113][31:0] = 32'd2830910537;
        ram[113][63:32] = 32'd2663013181;
        ram[113][95:64] = 32'd2238196546;
        ram[113][127:96] = 32'd3799628466;
        ram[114][31:0] = 32'd1297742875;
        ram[114][63:32] = 32'd2700525639;
        ram[114][95:64] = 32'd1845881788;
        ram[114][127:96] = 32'd582707416;
        ram[115][31:0] = 32'd3277373807;
        ram[115][63:32] = 32'd2115382646;
        ram[115][95:64] = 32'd3445572193;
        ram[115][127:96] = 32'd3340434727;
        ram[116][31:0] = 32'd1701612275;
        ram[116][63:32] = 32'd2952264133;
        ram[116][95:64] = 32'd2807963646;
        ram[116][127:96] = 32'd962725890;
        ram[117][31:0] = 32'd1954085459;
        ram[117][63:32] = 32'd1191579314;
        ram[117][95:64] = 32'd1183712898;
        ram[117][127:96] = 32'd987847086;
        ram[118][31:0] = 32'd2446660300;
        ram[118][63:32] = 32'd2376303146;
        ram[118][95:64] = 32'd107046119;
        ram[118][127:96] = 32'd1588844006;
        ram[119][31:0] = 32'd3484692570;
        ram[119][63:32] = 32'd702771066;
        ram[119][95:64] = 32'd3853924173;
        ram[119][127:96] = 32'd2750306313;
        ram[120][31:0] = 32'd1372344996;
        ram[120][63:32] = 32'd3284726031;
        ram[120][95:64] = 32'd2222178533;
        ram[120][127:96] = 32'd3017205182;
        ram[121][31:0] = 32'd1185966804;
        ram[121][63:32] = 32'd2138632015;
        ram[121][95:64] = 32'd2334539005;
        ram[121][127:96] = 32'd3597154848;
        ram[122][31:0] = 32'd1586990541;
        ram[122][63:32] = 32'd1052556506;
        ram[122][95:64] = 32'd541064026;
        ram[122][127:96] = 32'd2450647386;
        ram[123][31:0] = 32'd1030940358;
        ram[123][63:32] = 32'd1126176295;
        ram[123][95:64] = 32'd1405101754;
        ram[123][127:96] = 32'd1266991624;
        ram[124][31:0] = 32'd1858394599;
        ram[124][63:32] = 32'd2724175409;
        ram[124][95:64] = 32'd864413957;
        ram[124][127:96] = 32'd2620324755;
        ram[125][31:0] = 32'd1324133867;
        ram[125][63:32] = 32'd2750530624;
        ram[125][95:64] = 32'd2608397649;
        ram[125][127:96] = 32'd170019188;
        ram[126][31:0] = 32'd602751838;
        ram[126][63:32] = 32'd1706057765;
        ram[126][95:64] = 32'd846958545;
        ram[126][127:96] = 32'd640223175;
        ram[127][31:0] = 32'd1173294512;
        ram[127][63:32] = 32'd2952120113;
        ram[127][95:64] = 32'd154773377;
        ram[127][127:96] = 32'd1869058888;
        ram[128][31:0] = 32'd283576485;
        ram[128][63:32] = 32'd3832833658;
        ram[128][95:64] = 32'd1019661124;
        ram[128][127:96] = 32'd4175963926;
        ram[129][31:0] = 32'd2970200192;
        ram[129][63:32] = 32'd809825092;
        ram[129][95:64] = 32'd4077101732;
        ram[129][127:96] = 32'd1594848324;
        ram[130][31:0] = 32'd2499178703;
        ram[130][63:32] = 32'd4090293443;
        ram[130][95:64] = 32'd2119484876;
        ram[130][127:96] = 32'd2084861691;
        ram[131][31:0] = 32'd4169713201;
        ram[131][63:32] = 32'd2372613957;
        ram[131][95:64] = 32'd3622896168;
        ram[131][127:96] = 32'd1738182943;
        ram[132][31:0] = 32'd3364509141;
        ram[132][63:32] = 32'd2040683980;
        ram[132][95:64] = 32'd1199134247;
        ram[132][127:96] = 32'd3623927974;
        ram[133][31:0] = 32'd1098075619;
        ram[133][63:32] = 32'd3475139587;
        ram[133][95:64] = 32'd627486554;
        ram[133][127:96] = 32'd2501250615;
        ram[134][31:0] = 32'd4241396361;
        ram[134][63:32] = 32'd1845215902;
        ram[134][95:64] = 32'd2288013246;
        ram[134][127:96] = 32'd2749828337;
        ram[135][31:0] = 32'd30470061;
        ram[135][63:32] = 32'd2310349212;
        ram[135][95:64] = 32'd2967622748;
        ram[135][127:96] = 32'd1393884690;
        ram[136][31:0] = 32'd3477380391;
        ram[136][63:32] = 32'd87100184;
        ram[136][95:64] = 32'd1440277870;
        ram[136][127:96] = 32'd3210837133;
        ram[137][31:0] = 32'd1180199925;
        ram[137][63:32] = 32'd3421270430;
        ram[137][95:64] = 32'd2009710279;
        ram[137][127:96] = 32'd318746959;
        ram[138][31:0] = 32'd1846493572;
        ram[138][63:32] = 32'd298968730;
        ram[138][95:64] = 32'd3262924390;
        ram[138][127:96] = 32'd449821878;
        ram[139][31:0] = 32'd2994603037;
        ram[139][63:32] = 32'd2415573794;
        ram[139][95:64] = 32'd3010760443;
        ram[139][127:96] = 32'd455792188;
        ram[140][31:0] = 32'd4054210877;
        ram[140][63:32] = 32'd1362019700;
        ram[140][95:64] = 32'd286708441;
        ram[140][127:96] = 32'd38688635;
        ram[141][31:0] = 32'd2631069284;
        ram[141][63:32] = 32'd3264791009;
        ram[141][95:64] = 32'd3270728084;
        ram[141][127:96] = 32'd1469709198;
        ram[142][31:0] = 32'd352858729;
        ram[142][63:32] = 32'd1734513920;
        ram[142][95:64] = 32'd4085183514;
        ram[142][127:96] = 32'd2564920536;
        ram[143][31:0] = 32'd2320974549;
        ram[143][63:32] = 32'd1130181016;
        ram[143][95:64] = 32'd1311509596;
        ram[143][127:96] = 32'd1340627649;
        ram[144][31:0] = 32'd2352940238;
        ram[144][63:32] = 32'd861508937;
        ram[144][95:64] = 32'd3653426803;
        ram[144][127:96] = 32'd1094013198;
        ram[145][31:0] = 32'd1233267658;
        ram[145][63:32] = 32'd962066425;
        ram[145][95:64] = 32'd3179541911;
        ram[145][127:96] = 32'd2231704842;
        ram[146][31:0] = 32'd1490217735;
        ram[146][63:32] = 32'd1270660057;
        ram[146][95:64] = 32'd1844798620;
        ram[146][127:96] = 32'd3561949575;
        ram[147][31:0] = 32'd1893529001;
        ram[147][63:32] = 32'd1464251075;
        ram[147][95:64] = 32'd2083229337;
        ram[147][127:96] = 32'd3799185599;
        ram[148][31:0] = 32'd1467139886;
        ram[148][63:32] = 32'd704520665;
        ram[148][95:64] = 32'd499927349;
        ram[148][127:96] = 32'd2612499855;
        ram[149][31:0] = 32'd2164998835;
        ram[149][63:32] = 32'd4286678215;
        ram[149][95:64] = 32'd3698561184;
        ram[149][127:96] = 32'd2621666958;
        ram[150][31:0] = 32'd1153338480;
        ram[150][63:32] = 32'd647592843;
        ram[150][95:64] = 32'd1228005140;
        ram[150][127:96] = 32'd434815353;
        ram[151][31:0] = 32'd152904658;
        ram[151][63:32] = 32'd4068052147;
        ram[151][95:64] = 32'd906696308;
        ram[151][127:96] = 32'd2312933189;
        ram[152][31:0] = 32'd3635138265;
        ram[152][63:32] = 32'd1081248689;
        ram[152][95:64] = 32'd2988230185;
        ram[152][127:96] = 32'd701615759;
        ram[153][31:0] = 32'd2469017315;
        ram[153][63:32] = 32'd3646976116;
        ram[153][95:64] = 32'd2005415173;
        ram[153][127:96] = 32'd1197760716;
        ram[154][31:0] = 32'd1306428470;
        ram[154][63:32] = 32'd4082994306;
        ram[154][95:64] = 32'd902420674;
        ram[154][127:96] = 32'd2051461989;
        ram[155][31:0] = 32'd3343656720;
        ram[155][63:32] = 32'd723470077;
        ram[155][95:64] = 32'd2703610506;
        ram[155][127:96] = 32'd2813751329;
        ram[156][31:0] = 32'd2812841878;
        ram[156][63:32] = 32'd2462103418;
        ram[156][95:64] = 32'd2876902535;
        ram[156][127:96] = 32'd2689636519;
        ram[157][31:0] = 32'd2469942537;
        ram[157][63:32] = 32'd334721742;
        ram[157][95:64] = 32'd3572526873;
        ram[157][127:96] = 32'd842599967;
        ram[158][31:0] = 32'd3201343516;
        ram[158][63:32] = 32'd1874676766;
        ram[158][95:64] = 32'd954992338;
        ram[158][127:96] = 32'd2466428267;
        ram[159][31:0] = 32'd4218479966;
        ram[159][63:32] = 32'd1621771232;
        ram[159][95:64] = 32'd881995127;
        ram[159][127:96] = 32'd1193599707;
        ram[160][31:0] = 32'd1559299331;
        ram[160][63:32] = 32'd2087204287;
        ram[160][95:64] = 32'd1185904961;
        ram[160][127:96] = 32'd4156477301;
        ram[161][31:0] = 32'd3175733827;
        ram[161][63:32] = 32'd2042867590;
        ram[161][95:64] = 32'd4118931118;
        ram[161][127:96] = 32'd3927182985;
        ram[162][31:0] = 32'd3673972943;
        ram[162][63:32] = 32'd2151483163;
        ram[162][95:64] = 32'd1479657925;
        ram[162][127:96] = 32'd2006915388;
        ram[163][31:0] = 32'd3998291136;
        ram[163][63:32] = 32'd968066838;
        ram[163][95:64] = 32'd965599957;
        ram[163][127:96] = 32'd1564587862;
        ram[164][31:0] = 32'd1587342591;
        ram[164][63:32] = 32'd2971496127;
        ram[164][95:64] = 32'd501484569;
        ram[164][127:96] = 32'd4171986551;
        ram[165][31:0] = 32'd3089242911;
        ram[165][63:32] = 32'd507482648;
        ram[165][95:64] = 32'd267636255;
        ram[165][127:96] = 32'd2975358863;
        ram[166][31:0] = 32'd3762895607;
        ram[166][63:32] = 32'd1007391439;
        ram[166][95:64] = 32'd3229102402;
        ram[166][127:96] = 32'd243584986;
        ram[167][31:0] = 32'd4214335755;
        ram[167][63:32] = 32'd879311410;
        ram[167][95:64] = 32'd2700477505;
        ram[167][127:96] = 32'd3754236325;
        ram[168][31:0] = 32'd3988690396;
        ram[168][63:32] = 32'd1252547980;
        ram[168][95:64] = 32'd993674477;
        ram[168][127:96] = 32'd951086958;
        ram[169][31:0] = 32'd2458873297;
        ram[169][63:32] = 32'd3780631796;
        ram[169][95:64] = 32'd2431021203;
        ram[169][127:96] = 32'd2933532045;
        ram[170][31:0] = 32'd1881433713;
        ram[170][63:32] = 32'd1760731286;
        ram[170][95:64] = 32'd3793810237;
        ram[170][127:96] = 32'd1205808495;
        ram[171][31:0] = 32'd4251338616;
        ram[171][63:32] = 32'd1848469040;
        ram[171][95:64] = 32'd3756581141;
        ram[171][127:96] = 32'd258286431;
        ram[172][31:0] = 32'd3658468012;
        ram[172][63:32] = 32'd1050422211;
        ram[172][95:64] = 32'd2572045592;
        ram[172][127:96] = 32'd1533424138;
        ram[173][31:0] = 32'd1185532734;
        ram[173][63:32] = 32'd1966776275;
        ram[173][95:64] = 32'd3428477096;
        ram[173][127:96] = 32'd2233471613;
        ram[174][31:0] = 32'd510585055;
        ram[174][63:32] = 32'd241466137;
        ram[174][95:64] = 32'd1941058159;
        ram[174][127:96] = 32'd2964207096;
        ram[175][31:0] = 32'd4290278596;
        ram[175][63:32] = 32'd3363580375;
        ram[175][95:64] = 32'd1769260887;
        ram[175][127:96] = 32'd892604545;
        ram[176][31:0] = 32'd2931391489;
        ram[176][63:32] = 32'd2046342139;
        ram[176][95:64] = 32'd1271505191;
        ram[176][127:96] = 32'd986566342;
        ram[177][31:0] = 32'd2576467063;
        ram[177][63:32] = 32'd83794451;
        ram[177][95:64] = 32'd2751230606;
        ram[177][127:96] = 32'd3928838089;
        ram[178][31:0] = 32'd2682563090;
        ram[178][63:32] = 32'd3261845956;
        ram[178][95:64] = 32'd4226705526;
        ram[178][127:96] = 32'd3264214500;
        ram[179][31:0] = 32'd3183387761;
        ram[179][63:32] = 32'd3532130073;
        ram[179][95:64] = 32'd2494614555;
        ram[179][127:96] = 32'd2722927766;
        ram[180][31:0] = 32'd2104937406;
        ram[180][63:32] = 32'd2025627376;
        ram[180][95:64] = 32'd3889326331;
        ram[180][127:96] = 32'd3748128516;
        ram[181][31:0] = 32'd1310629757;
        ram[181][63:32] = 32'd3136553366;
        ram[181][95:64] = 32'd1207862729;
        ram[181][127:96] = 32'd1005793312;
        ram[182][31:0] = 32'd2860904189;
        ram[182][63:32] = 32'd2983101154;
        ram[182][95:64] = 32'd3958101048;
        ram[182][127:96] = 32'd1353510671;
        ram[183][31:0] = 32'd848268891;
        ram[183][63:32] = 32'd1312293725;
        ram[183][95:64] = 32'd3494088879;
        ram[183][127:96] = 32'd567958459;
        ram[184][31:0] = 32'd967452695;
        ram[184][63:32] = 32'd276361428;
        ram[184][95:64] = 32'd791004845;
        ram[184][127:96] = 32'd3426545964;
        ram[185][31:0] = 32'd574474385;
        ram[185][63:32] = 32'd1810153704;
        ram[185][95:64] = 32'd2878401245;
        ram[185][127:96] = 32'd292010483;
        ram[186][31:0] = 32'd230455895;
        ram[186][63:32] = 32'd3435630877;
        ram[186][95:64] = 32'd3185922216;
        ram[186][127:96] = 32'd2859145874;
        ram[187][31:0] = 32'd3916469345;
        ram[187][63:32] = 32'd1248251572;
        ram[187][95:64] = 32'd282558174;
        ram[187][127:96] = 32'd3419461017;
        ram[188][31:0] = 32'd467983000;
        ram[188][63:32] = 32'd3215843439;
        ram[188][95:64] = 32'd2930249500;
        ram[188][127:96] = 32'd997232407;
        ram[189][31:0] = 32'd1081173468;
        ram[189][63:32] = 32'd2619751839;
        ram[189][95:64] = 32'd1230763844;
        ram[189][127:96] = 32'd1446998705;
        ram[190][31:0] = 32'd3811051108;
        ram[190][63:32] = 32'd3770741534;
        ram[190][95:64] = 32'd3993692466;
        ram[190][127:96] = 32'd930239523;
        ram[191][31:0] = 32'd2449701785;
        ram[191][63:32] = 32'd3541645589;
        ram[191][95:64] = 32'd910969802;
        ram[191][127:96] = 32'd2089824228;
        ram[192][31:0] = 32'd4228114320;
        ram[192][63:32] = 32'd3880414256;
        ram[192][95:64] = 32'd317508578;
        ram[192][127:96] = 32'd2119250569;
        ram[193][31:0] = 32'd1620593328;
        ram[193][63:32] = 32'd256807720;
        ram[193][95:64] = 32'd9534195;
        ram[193][127:96] = 32'd4171009354;
        ram[194][31:0] = 32'd3596983855;
        ram[194][63:32] = 32'd3617657151;
        ram[194][95:64] = 32'd1257411684;
        ram[194][127:96] = 32'd312513893;
        ram[195][31:0] = 32'd1167957788;
        ram[195][63:32] = 32'd3802541709;
        ram[195][95:64] = 32'd3995135572;
        ram[195][127:96] = 32'd973592663;
        ram[196][31:0] = 32'd10366515;
        ram[196][63:32] = 32'd3660035070;
        ram[196][95:64] = 32'd3459446628;
        ram[196][127:96] = 32'd3341782422;
        ram[197][31:0] = 32'd1105670773;
        ram[197][63:32] = 32'd911008138;
        ram[197][95:64] = 32'd1470099950;
        ram[197][127:96] = 32'd785259291;
        ram[198][31:0] = 32'd626252886;
        ram[198][63:32] = 32'd1321282978;
        ram[198][95:64] = 32'd4231216897;
        ram[198][127:96] = 32'd1922871569;
        ram[199][31:0] = 32'd2646907564;
        ram[199][63:32] = 32'd99933581;
        ram[199][95:64] = 32'd3837150160;
        ram[199][127:96] = 32'd3441245320;
        ram[200][31:0] = 32'd3100164281;
        ram[200][63:32] = 32'd1686375627;
        ram[200][95:64] = 32'd4239473607;
        ram[200][127:96] = 32'd4046978904;
        ram[201][31:0] = 32'd1315671584;
        ram[201][63:32] = 32'd3455870968;
        ram[201][95:64] = 32'd1359101487;
        ram[201][127:96] = 32'd540490609;
        ram[202][31:0] = 32'd4179863201;
        ram[202][63:32] = 32'd4112399394;
        ram[202][95:64] = 32'd3925951955;
        ram[202][127:96] = 32'd4155520991;
        ram[203][31:0] = 32'd3444397451;
        ram[203][63:32] = 32'd3209556232;
        ram[203][95:64] = 32'd3061961020;
        ram[203][127:96] = 32'd99083937;
        ram[204][31:0] = 32'd3371550778;
        ram[204][63:32] = 32'd3864354102;
        ram[204][95:64] = 32'd3123056303;
        ram[204][127:96] = 32'd2697333757;
        ram[205][31:0] = 32'd1650346404;
        ram[205][63:32] = 32'd971615072;
        ram[205][95:64] = 32'd2907326481;
        ram[205][127:96] = 32'd532265002;
        ram[206][31:0] = 32'd3204893334;
        ram[206][63:32] = 32'd2120594327;
        ram[206][95:64] = 32'd2805664193;
        ram[206][127:96] = 32'd1406447338;
        ram[207][31:0] = 32'd1271401654;
        ram[207][63:32] = 32'd3795551779;
        ram[207][95:64] = 32'd72105947;
        ram[207][127:96] = 32'd2426107502;
        ram[208][31:0] = 32'd4001181699;
        ram[208][63:32] = 32'd1217572098;
        ram[208][95:64] = 32'd4233557749;
        ram[208][127:96] = 32'd3366828491;
        ram[209][31:0] = 32'd4021549176;
        ram[209][63:32] = 32'd1959645325;
        ram[209][95:64] = 32'd3573850885;
        ram[209][127:96] = 32'd1323733114;
        ram[210][31:0] = 32'd1623547379;
        ram[210][63:32] = 32'd729735648;
        ram[210][95:64] = 32'd3905935845;
        ram[210][127:96] = 32'd64812169;
        ram[211][31:0] = 32'd1905889562;
        ram[211][63:32] = 32'd3605691528;
        ram[211][95:64] = 32'd3157279990;
        ram[211][127:96] = 32'd4178636307;
        ram[212][31:0] = 32'd1091101872;
        ram[212][63:32] = 32'd2875037109;
        ram[212][95:64] = 32'd1086596891;
        ram[212][127:96] = 32'd30109657;
        ram[213][31:0] = 32'd201249939;
        ram[213][63:32] = 32'd1375294070;
        ram[213][95:64] = 32'd3733979249;
        ram[213][127:96] = 32'd3155227187;
        ram[214][31:0] = 32'd3338308047;
        ram[214][63:32] = 32'd904680371;
        ram[214][95:64] = 32'd3668307118;
        ram[214][127:96] = 32'd790427723;
        ram[215][31:0] = 32'd2040878775;
        ram[215][63:32] = 32'd2853075293;
        ram[215][95:64] = 32'd3234096972;
        ram[215][127:96] = 32'd983979571;
        ram[216][31:0] = 32'd2537001022;
        ram[216][63:32] = 32'd3049915918;
        ram[216][95:64] = 32'd2528451676;
        ram[216][127:96] = 32'd4195620311;
        ram[217][31:0] = 32'd749785393;
        ram[217][63:32] = 32'd3921532732;
        ram[217][95:64] = 32'd1773147721;
        ram[217][127:96] = 32'd3229558777;
        ram[218][31:0] = 32'd1918914483;
        ram[218][63:32] = 32'd1520019581;
        ram[218][95:64] = 32'd2978499719;
        ram[218][127:96] = 32'd1778218794;
        ram[219][31:0] = 32'd3812382912;
        ram[219][63:32] = 32'd2926156055;
        ram[219][95:64] = 32'd1560394632;
        ram[219][127:96] = 32'd4177420437;
        ram[220][31:0] = 32'd1391719360;
        ram[220][63:32] = 32'd1878584955;
        ram[220][95:64] = 32'd2047159171;
        ram[220][127:96] = 32'd3827280495;
        ram[221][31:0] = 32'd700616692;
        ram[221][63:32] = 32'd3458389258;
        ram[221][95:64] = 32'd3642098538;
        ram[221][127:96] = 32'd2507313658;
        ram[222][31:0] = 32'd397640837;
        ram[222][63:32] = 32'd1528309135;
        ram[222][95:64] = 32'd42358296;
        ram[222][127:96] = 32'd1369333498;
        ram[223][31:0] = 32'd3751642818;
        ram[223][63:32] = 32'd2422299734;
        ram[223][95:64] = 32'd585438621;
        ram[223][127:96] = 32'd3072952231;
        ram[224][31:0] = 32'd819431204;
        ram[224][63:32] = 32'd268761716;
        ram[224][95:64] = 32'd2940907252;
        ram[224][127:96] = 32'd4140880084;
        ram[225][31:0] = 32'd3274897863;
        ram[225][63:32] = 32'd179229824;
        ram[225][95:64] = 32'd3561446271;
        ram[225][127:96] = 32'd486481265;
        ram[226][31:0] = 32'd299855562;
        ram[226][63:32] = 32'd1328078859;
        ram[226][95:64] = 32'd487641621;
        ram[226][127:96] = 32'd1829404985;
        ram[227][31:0] = 32'd3676688916;
        ram[227][63:32] = 32'd3145412611;
        ram[227][95:64] = 32'd518895518;
        ram[227][127:96] = 32'd806648968;
        ram[228][31:0] = 32'd3690236031;
        ram[228][63:32] = 32'd858191111;
        ram[228][95:64] = 32'd4191420171;
        ram[228][127:96] = 32'd2854654772;
        ram[229][31:0] = 32'd936149391;
        ram[229][63:32] = 32'd3442910521;
        ram[229][95:64] = 32'd3381071146;
        ram[229][127:96] = 32'd632463510;
        ram[230][31:0] = 32'd1241003816;
        ram[230][63:32] = 32'd3835640528;
        ram[230][95:64] = 32'd2267903388;
        ram[230][127:96] = 32'd3334114139;
        ram[231][31:0] = 32'd2084629605;
        ram[231][63:32] = 32'd2610089944;
        ram[231][95:64] = 32'd1323017946;
        ram[231][127:96] = 32'd425505923;
        ram[232][31:0] = 32'd1778724627;
        ram[232][63:32] = 32'd2967891672;
        ram[232][95:64] = 32'd1564872363;
        ram[232][127:96] = 32'd4191689811;
        ram[233][31:0] = 32'd572260113;
        ram[233][63:32] = 32'd1769109334;
        ram[233][95:64] = 32'd1484061370;
        ram[233][127:96] = 32'd2013495484;
        ram[234][31:0] = 32'd607348316;
        ram[234][63:32] = 32'd625389764;
        ram[234][95:64] = 32'd2087976953;
        ram[234][127:96] = 32'd2971125663;
        ram[235][31:0] = 32'd3211187226;
        ram[235][63:32] = 32'd1873325343;
        ram[235][95:64] = 32'd3185997769;
        ram[235][127:96] = 32'd1653503808;
        ram[236][31:0] = 32'd1934668787;
        ram[236][63:32] = 32'd1578395060;
        ram[236][95:64] = 32'd1984305920;
        ram[236][127:96] = 32'd2267174355;
        ram[237][31:0] = 32'd292043820;
        ram[237][63:32] = 32'd1182899197;
        ram[237][95:64] = 32'd2459752245;
        ram[237][127:96] = 32'd3631193825;
        ram[238][31:0] = 32'd1791314849;
        ram[238][63:32] = 32'd2693867941;
        ram[238][95:64] = 32'd613951372;
        ram[238][127:96] = 32'd905894982;
        ram[239][31:0] = 32'd90020364;
        ram[239][63:32] = 32'd2991872276;
        ram[239][95:64] = 32'd3447221745;
        ram[239][127:96] = 32'd1132988677;
        ram[240][31:0] = 32'd307012169;
        ram[240][63:32] = 32'd762603117;
        ram[240][95:64] = 32'd2765447673;
        ram[240][127:96] = 32'd313403234;
        ram[241][31:0] = 32'd3129425578;
        ram[241][63:32] = 32'd628646139;
        ram[241][95:64] = 32'd2560894838;
        ram[241][127:96] = 32'd2075372781;
        ram[242][31:0] = 32'd3571431660;
        ram[242][63:32] = 32'd682498780;
        ram[242][95:64] = 32'd4208904194;
        ram[242][127:96] = 32'd1365898262;
        ram[243][31:0] = 32'd1158453115;
        ram[243][63:32] = 32'd3512163126;
        ram[243][95:64] = 32'd1819208149;
        ram[243][127:96] = 32'd900993035;
        ram[244][31:0] = 32'd888555328;
        ram[244][63:32] = 32'd871000283;
        ram[244][95:64] = 32'd1143928461;
        ram[244][127:96] = 32'd3552257411;
        ram[245][31:0] = 32'd1860707669;
        ram[245][63:32] = 32'd3490086291;
        ram[245][95:64] = 32'd327157360;
        ram[245][127:96] = 32'd3859842153;
        ram[246][31:0] = 32'd447706912;
        ram[246][63:32] = 32'd3871310064;
        ram[246][95:64] = 32'd2041805604;
        ram[246][127:96] = 32'd730636411;
        ram[247][31:0] = 32'd1189533474;
        ram[247][63:32] = 32'd3261557463;
        ram[247][95:64] = 32'd431413773;
        ram[247][127:96] = 32'd961558183;
        ram[248][31:0] = 32'd1625093277;
        ram[248][63:32] = 32'd1150199168;
        ram[248][95:64] = 32'd3736541262;
        ram[248][127:96] = 32'd1594198084;
        ram[249][31:0] = 32'd103670533;
        ram[249][63:32] = 32'd2851191842;
        ram[249][95:64] = 32'd856833474;
        ram[249][127:96] = 32'd811944595;
        ram[250][31:0] = 32'd2148363208;
        ram[250][63:32] = 32'd3133226956;
        ram[250][95:64] = 32'd1816079453;
        ram[250][127:96] = 32'd3753928122;
        ram[251][31:0] = 32'd4090172265;
        ram[251][63:32] = 32'd1735952530;
        ram[251][95:64] = 32'd1873145601;
        ram[251][127:96] = 32'd635148783;
        ram[252][31:0] = 32'd2350202510;
        ram[252][63:32] = 32'd3720685503;
        ram[252][95:64] = 32'd1146572673;
        ram[252][127:96] = 32'd1935275313;
        ram[253][31:0] = 32'd128963949;
        ram[253][63:32] = 32'd3119782812;
        ram[253][95:64] = 32'd2391167737;
        ram[253][127:96] = 32'd8870532;
        ram[254][31:0] = 32'd2828332147;
        ram[254][63:32] = 32'd3197795730;
        ram[254][95:64] = 32'd2750972131;
        ram[254][127:96] = 32'd754054502;
        ram[255][31:0] = 32'd1322191517;
        ram[255][63:32] = 32'd46789532;
        ram[255][95:64] = 32'd2746665182;
        ram[255][127:96] = 32'd4086440552;

    end
    always @(posedge clk) begin
        addr_r <= raddr;
        if(we) ram[waddr] <= din;
    end
    assign dout = ram[addr_r]; 

endmodule

//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/03/31 14:48:12
// Design Name: 
// Module Name: PC
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module PC (
    input                   [ 0 : 0]            clk,
    input                   [ 0 : 0]            rst,
    input                   [ 0 : 0]            en,
    input                   [ 0 : 0]            flush,
    input                   [ 0 : 0]            stall,
    input                   [31 : 0]            npc,
    output      reg         [31 : 0]            pc
);

always @(posedge clk) begin
    if(rst)
        pc<=32'H00400000;
    else if (en) begin
        if (flush) begin
            pc<=npc;
        end
        else if (!stall) begin
            pc<=npc;
        end
    end
end

endmodule


/*
本文件是一个测试文件，用于测试cache模块
工作原理是模仿CPU的读写请求，对cache进行读写操作
将Cache返回的数据与预先数据进行比较，如果一致则测试通过
*/
`timescale 1ns/1ps
module cache_tb();

    //测试参数
    parameter READ_NUM = 2000;  // 测试次数 这里设置为2000次读，1000次写
    parameter WRITE_NUM = 1000;  
    //模块参数
    parameter INDEX_WIDTH       = 2;   // Cache索引位宽 2^3=8行
    parameter LINE_OFFSET_WIDTH = 2;   // 行偏移位宽，决定了一行的宽度 2^2=4字
    parameter SPACE_OFFSET      = 2;   // 一个地址空间占1个字节，因此一个字需要4个地址空间，由于假设为整字读取，处理地址的时候可以默认后两位为0
    parameter MEM_ADDR_WIDTH    = 10;   // 为了简化，这里假设内存地址宽度为10位（CPU请求地址仍然是32位，只不过我们这里简化处理，截断了高位） 
    parameter WAY_NUM           = 2;   // Cache N路组相联(N=1的时候是直接映射)
    parameter REPLACE_POLICY    = 0;   // 替换策略 0：LRU 1：FIFO 2：伪随机

    // 变化的信号 CPU发出
    reg clk=1;
    reg rstn=1;
    reg stat=0;
    // 等rstn信号稳定后 clk信号才开始翻转
    initial begin
        #1 rstn = 0;
        #1 rstn = 1;
        stat = 1;
    end
    always  #1 clk = ~clk;

    wire [31:0] addr;
    wire r_req;
    wire w_req;
    wire [31:0] w_data;

    // 导线
    wire [31:0] r_data;
    wire miss;
    wire mem_r;
    wire mem_w;
    wire [31:0] mem_addr;
    wire [127:0] mem_w_data;
    wire [127:0] mem_r_data;
    wire mem_ready;

    // 用于测试的信号
    reg [MEM_ADDR_WIDTH-1:0] test_addr[0:READ_NUM+WRITE_NUM-1];  // 用于存储测试地址
    reg [32:0] test_data[0:READ_NUM+WRITE_NUM-1];  // 用于存储测试数据 最高位用于标记是否写入 0：读 1：写
    reg [31:0] test_cnt=0;  // 用于计数，每次读写操作后加1
    reg diff=0;  // 用于标记是否有不一致的数据

    // 用于对比的提交，当前cache应该给出的数据
    wire op;
    wire[31:0] data;
    assign op = test_data[test_cnt-1][32];
    assign data = test_data[test_cnt-1][31:0];
    
    // 状态机
    assign addr = test_addr[test_cnt]<<SPACE_OFFSET;
    assign r_req = test_data[test_cnt][32] == 0 ? 1 : 0;
    assign w_req = test_data[test_cnt][32] == 1 ? 1 : 0;
    assign w_data = test_data[test_cnt][31:0];
    always @(posedge clk) begin
        if (!miss && (test_cnt < READ_NUM+WRITE_NUM) && stat) begin
            if (test_data[test_cnt-1][32] == 0) begin  // 读
                if (r_data != test_data[test_cnt-1][31:0]) begin
                    $display("Read error at %d, expect %h, get %h", test_cnt, test_data[test_cnt-1][31:0], r_data);
                    diff = 1;
                end
            end
            test_cnt <= test_cnt + 1;
        end
    end

    // 例化cache
    cache #(
        .INDEX_WIDTH(INDEX_WIDTH),
        .LINE_OFFSET_WIDTH(LINE_OFFSET_WIDTH),
        .SPACE_OFFSET(SPACE_OFFSET),
        .WAY_NUM(WAY_NUM),
        .REPLACE_POLICY(REPLACE_POLICY)
    ) cache_inst(
        .clk(clk),
        .rstn(rstn),
        .addr(addr),
        .r_req(r_req),
        .w_req(w_req),
        .w_data(w_data),
        .r_data(r_data),
        .miss(miss),
        .mem_r(mem_r),
        .mem_w(mem_w),
        .mem_addr(mem_addr),
        .mem_w_data(mem_w_data),
        .mem_r_data(mem_r_data),
        .mem_ready(mem_ready)
    );

    // 内存
    mem #(
        .INDEX_WIDTH(INDEX_WIDTH),
        .LINE_OFFSET_WIDTH(LINE_OFFSET_WIDTH),
        .SPACE_OFFSET(SPACE_OFFSET),
        .MEM_ADDR_WIDTH(MEM_ADDR_WIDTH-LINE_OFFSET_WIDTH),
        .WAY_NUM(WAY_NUM)
    ) mem_inst(
        .clk(clk),
        .rstn(rstn),
        .mem_r(mem_r),
        .mem_w(mem_w),
        .mem_addr(mem_addr),
        .mem_w_data(mem_w_data),
        .mem_r_data(mem_r_data),
        .mem_ready(mem_ready)
    );

    // 初始化测试数据
    initial begin
        test_addr[0] = 960;
        test_data[0] = 33'd5729732664;
        test_addr[1] = 576;
        test_data[1] = 33'd2373603425;
        test_addr[2] = 810;
        test_data[2] = 33'd1557606680;
        test_addr[3] = 13;
        test_data[3] = 33'd1541123444;
        test_addr[4] = 358;
        test_data[4] = 33'd3979567529;
        test_addr[5] = 920;
        test_data[5] = 33'd3925196331;
        test_addr[6] = 307;
        test_data[6] = 33'd6852386940;
        test_addr[7] = 457;
        test_data[7] = 33'd5073763691;
        test_addr[8] = 221;
        test_data[8] = 33'd5015325859;
        test_addr[9] = 818;
        test_data[9] = 33'd2986767408;
        test_addr[10] = 822;
        test_data[10] = 33'd534736813;
        test_addr[11] = 1009;
        test_data[11] = 33'd2054454801;
        test_addr[12] = 905;
        test_data[12] = 33'd3362997925;
        test_addr[13] = 896;
        test_data[13] = 33'd7920708864;
        test_addr[14] = 558;
        test_data[14] = 33'd3650811963;
        test_addr[15] = 565;
        test_data[15] = 33'd7138605058;
        test_addr[16] = 184;
        test_data[16] = 33'd8135532124;
        test_addr[17] = 657;
        test_data[17] = 33'd3120162192;
        test_addr[18] = 631;
        test_data[18] = 33'd7920984454;
        test_addr[19] = 74;
        test_data[19] = 33'd3405503829;
        test_addr[20] = 720;
        test_data[20] = 33'd2954885626;
        test_addr[21] = 164;
        test_data[21] = 33'd6072879824;
        test_addr[22] = 379;
        test_data[22] = 33'd1897669063;
        test_addr[23] = 713;
        test_data[23] = 33'd333588719;
        test_addr[24] = 961;
        test_data[24] = 33'd2071565022;
        test_addr[25] = 461;
        test_data[25] = 33'd4299739377;
        test_addr[26] = 858;
        test_data[26] = 33'd2562306931;
        test_addr[27] = 856;
        test_data[27] = 33'd975862316;
        test_addr[28] = 824;
        test_data[28] = 33'd3205965066;
        test_addr[29] = 683;
        test_data[29] = 33'd3865309988;
        test_addr[30] = 0;
        test_data[30] = 33'd7509293195;
        test_addr[31] = 812;
        test_data[31] = 33'd2625492882;
        test_addr[32] = 467;
        test_data[32] = 33'd8128350892;
        test_addr[33] = 461;
        test_data[33] = 33'd4772081;
        test_addr[34] = 754;
        test_data[34] = 33'd5526759199;
        test_addr[35] = 249;
        test_data[35] = 33'd3978129519;
        test_addr[36] = 273;
        test_data[36] = 33'd56693191;
        test_addr[37] = 379;
        test_data[37] = 33'd7543914694;
        test_addr[38] = 304;
        test_data[38] = 33'd3014575534;
        test_addr[39] = 423;
        test_data[39] = 33'd5858825227;
        test_addr[40] = 918;
        test_data[40] = 33'd2681524291;
        test_addr[41] = 727;
        test_data[41] = 33'd2717525231;
        test_addr[42] = 1001;
        test_data[42] = 33'd6113713893;
        test_addr[43] = 513;
        test_data[43] = 33'd8012642441;
        test_addr[44] = 353;
        test_data[44] = 33'd3399552858;
        test_addr[45] = 919;
        test_data[45] = 33'd4642040004;
        test_addr[46] = 826;
        test_data[46] = 33'd4985112467;
        test_addr[47] = 616;
        test_data[47] = 33'd2000952156;
        test_addr[48] = 658;
        test_data[48] = 33'd5527266926;
        test_addr[49] = 377;
        test_data[49] = 33'd6665831953;
        test_addr[50] = 479;
        test_data[50] = 33'd3763673002;
        test_addr[51] = 930;
        test_data[51] = 33'd890973601;
        test_addr[52] = 523;
        test_data[52] = 33'd4872652897;
        test_addr[53] = 556;
        test_data[53] = 33'd2629206974;
        test_addr[54] = 508;
        test_data[54] = 33'd2569124247;
        test_addr[55] = 608;
        test_data[55] = 33'd7676707290;
        test_addr[56] = 141;
        test_data[56] = 33'd324907900;
        test_addr[57] = 989;
        test_data[57] = 33'd6581277516;
        test_addr[58] = 591;
        test_data[58] = 33'd4087477473;
        test_addr[59] = 276;
        test_data[59] = 33'd6989463839;
        test_addr[60] = 95;
        test_data[60] = 33'd8261569972;
        test_addr[61] = 154;
        test_data[61] = 33'd1881539630;
        test_addr[62] = 943;
        test_data[62] = 33'd6778659248;
        test_addr[63] = 29;
        test_data[63] = 33'd1848244721;
        test_addr[64] = 18;
        test_data[64] = 33'd4718483358;
        test_addr[65] = 2;
        test_data[65] = 33'd3771999802;
        test_addr[66] = 361;
        test_data[66] = 33'd5849023877;
        test_addr[67] = 615;
        test_data[67] = 33'd2136755942;
        test_addr[68] = 2;
        test_data[68] = 33'd3771999802;
        test_addr[69] = 865;
        test_data[69] = 33'd1605398418;
        test_addr[70] = 421;
        test_data[70] = 33'd2522318236;
        test_addr[71] = 503;
        test_data[71] = 33'd2825090233;
        test_addr[72] = 432;
        test_data[72] = 33'd926426471;
        test_addr[73] = 542;
        test_data[73] = 33'd6729107974;
        test_addr[74] = 80;
        test_data[74] = 33'd818068638;
        test_addr[75] = 176;
        test_data[75] = 33'd2275341057;
        test_addr[76] = 839;
        test_data[76] = 33'd5004566380;
        test_addr[77] = 728;
        test_data[77] = 33'd128590783;
        test_addr[78] = 508;
        test_data[78] = 33'd2569124247;
        test_addr[79] = 509;
        test_data[79] = 33'd1404134308;
        test_addr[80] = 633;
        test_data[80] = 33'd3083058234;
        test_addr[81] = 960;
        test_data[81] = 33'd1434765368;
        test_addr[82] = 286;
        test_data[82] = 33'd2360048588;
        test_addr[83] = 158;
        test_data[83] = 33'd217812934;
        test_addr[84] = 28;
        test_data[84] = 33'd1087055728;
        test_addr[85] = 940;
        test_data[85] = 33'd2787861430;
        test_addr[86] = 830;
        test_data[86] = 33'd2069122430;
        test_addr[87] = 129;
        test_data[87] = 33'd6177050060;
        test_addr[88] = 417;
        test_data[88] = 33'd6563850865;
        test_addr[89] = 897;
        test_data[89] = 33'd4367054241;
        test_addr[90] = 398;
        test_data[90] = 33'd1175204693;
        test_addr[91] = 408;
        test_data[91] = 33'd5425803462;
        test_addr[92] = 165;
        test_data[92] = 33'd106644142;
        test_addr[93] = 131;
        test_data[93] = 33'd5108247865;
        test_addr[94] = 375;
        test_data[94] = 33'd1408822660;
        test_addr[95] = 559;
        test_data[95] = 33'd3112428785;
        test_addr[96] = 6;
        test_data[96] = 33'd1280683540;
        test_addr[97] = 525;
        test_data[97] = 33'd4721499492;
        test_addr[98] = 420;
        test_data[98] = 33'd3817791626;
        test_addr[99] = 638;
        test_data[99] = 33'd7552127021;
        test_addr[100] = 483;
        test_data[100] = 33'd1178549137;
        test_addr[101] = 637;
        test_data[101] = 33'd1672692856;
        test_addr[102] = 179;
        test_data[102] = 33'd2011666985;
        test_addr[103] = 877;
        test_data[103] = 33'd5612476653;
        test_addr[104] = 547;
        test_data[104] = 33'd2109417922;
        test_addr[105] = 848;
        test_data[105] = 33'd415536288;
        test_addr[106] = 716;
        test_data[106] = 33'd5636059386;
        test_addr[107] = 81;
        test_data[107] = 33'd7686742519;
        test_addr[108] = 394;
        test_data[108] = 33'd496284610;
        test_addr[109] = 435;
        test_data[109] = 33'd3843532341;
        test_addr[110] = 929;
        test_data[110] = 33'd2947338001;
        test_addr[111] = 534;
        test_data[111] = 33'd1059137997;
        test_addr[112] = 654;
        test_data[112] = 33'd1773452330;
        test_addr[113] = 778;
        test_data[113] = 33'd3444963042;
        test_addr[114] = 430;
        test_data[114] = 33'd3947540049;
        test_addr[115] = 1016;
        test_data[115] = 33'd595270188;
        test_addr[116] = 966;
        test_data[116] = 33'd1835137690;
        test_addr[117] = 847;
        test_data[117] = 33'd196428976;
        test_addr[118] = 669;
        test_data[118] = 33'd2603095900;
        test_addr[119] = 130;
        test_data[119] = 33'd1268433295;
        test_addr[120] = 947;
        test_data[120] = 33'd965247601;
        test_addr[121] = 1023;
        test_data[121] = 33'd1969797033;
        test_addr[122] = 737;
        test_data[122] = 33'd3825165600;
        test_addr[123] = 583;
        test_data[123] = 33'd4069883337;
        test_addr[124] = 568;
        test_data[124] = 33'd2796273124;
        test_addr[125] = 228;
        test_data[125] = 33'd3498918036;
        test_addr[126] = 478;
        test_data[126] = 33'd4922267630;
        test_addr[127] = 577;
        test_data[127] = 33'd5126013402;
        test_addr[128] = 818;
        test_data[128] = 33'd2986767408;
        test_addr[129] = 381;
        test_data[129] = 33'd3910801142;
        test_addr[130] = 736;
        test_data[130] = 33'd65646729;
        test_addr[131] = 437;
        test_data[131] = 33'd3188866646;
        test_addr[132] = 65;
        test_data[132] = 33'd993562414;
        test_addr[133] = 710;
        test_data[133] = 33'd8543008649;
        test_addr[134] = 179;
        test_data[134] = 33'd7728460445;
        test_addr[135] = 139;
        test_data[135] = 33'd3677407724;
        test_addr[136] = 844;
        test_data[136] = 33'd1272998109;
        test_addr[137] = 1018;
        test_data[137] = 33'd3013633939;
        test_addr[138] = 183;
        test_data[138] = 33'd8006673390;
        test_addr[139] = 502;
        test_data[139] = 33'd7585331964;
        test_addr[140] = 956;
        test_data[140] = 33'd3817405510;
        test_addr[141] = 180;
        test_data[141] = 33'd4026446541;
        test_addr[142] = 251;
        test_data[142] = 33'd1773791810;
        test_addr[143] = 280;
        test_data[143] = 33'd761284035;
        test_addr[144] = 82;
        test_data[144] = 33'd1240469410;
        test_addr[145] = 459;
        test_data[145] = 33'd2890618210;
        test_addr[146] = 2;
        test_data[146] = 33'd3771999802;
        test_addr[147] = 740;
        test_data[147] = 33'd2129383015;
        test_addr[148] = 400;
        test_data[148] = 33'd545504374;
        test_addr[149] = 267;
        test_data[149] = 33'd7922293771;
        test_addr[150] = 173;
        test_data[150] = 33'd1456155483;
        test_addr[151] = 778;
        test_data[151] = 33'd3444963042;
        test_addr[152] = 897;
        test_data[152] = 33'd72086945;
        test_addr[153] = 632;
        test_data[153] = 33'd162213990;
        test_addr[154] = 10;
        test_data[154] = 33'd8380090129;
        test_addr[155] = 80;
        test_data[155] = 33'd818068638;
        test_addr[156] = 553;
        test_data[156] = 33'd4101269385;
        test_addr[157] = 824;
        test_data[157] = 33'd4606386530;
        test_addr[158] = 1015;
        test_data[158] = 33'd2062647632;
        test_addr[159] = 600;
        test_data[159] = 33'd1402039586;
        test_addr[160] = 906;
        test_data[160] = 33'd1312679890;
        test_addr[161] = 311;
        test_data[161] = 33'd7798885443;
        test_addr[162] = 925;
        test_data[162] = 33'd6078202650;
        test_addr[163] = 587;
        test_data[163] = 33'd702014159;
        test_addr[164] = 942;
        test_data[164] = 33'd8397752001;
        test_addr[165] = 308;
        test_data[165] = 33'd4977428107;
        test_addr[166] = 123;
        test_data[166] = 33'd3515538989;
        test_addr[167] = 627;
        test_data[167] = 33'd5605669470;
        test_addr[168] = 573;
        test_data[168] = 33'd3693245975;
        test_addr[169] = 741;
        test_data[169] = 33'd3239258243;
        test_addr[170] = 73;
        test_data[170] = 33'd5070048379;
        test_addr[171] = 343;
        test_data[171] = 33'd6767134447;
        test_addr[172] = 221;
        test_data[172] = 33'd720358563;
        test_addr[173] = 1009;
        test_data[173] = 33'd2054454801;
        test_addr[174] = 722;
        test_data[174] = 33'd4149935825;
        test_addr[175] = 846;
        test_data[175] = 33'd6358430626;
        test_addr[176] = 311;
        test_data[176] = 33'd3503918147;
        test_addr[177] = 163;
        test_data[177] = 33'd5935134857;
        test_addr[178] = 886;
        test_data[178] = 33'd4267669502;
        test_addr[179] = 221;
        test_data[179] = 33'd720358563;
        test_addr[180] = 198;
        test_data[180] = 33'd4018594710;
        test_addr[181] = 979;
        test_data[181] = 33'd5804725036;
        test_addr[182] = 49;
        test_data[182] = 33'd751512591;
        test_addr[183] = 780;
        test_data[183] = 33'd404411201;
        test_addr[184] = 940;
        test_data[184] = 33'd5053645011;
        test_addr[185] = 162;
        test_data[185] = 33'd1711500696;
        test_addr[186] = 595;
        test_data[186] = 33'd1438576721;
        test_addr[187] = 709;
        test_data[187] = 33'd1267071129;
        test_addr[188] = 459;
        test_data[188] = 33'd7102986280;
        test_addr[189] = 385;
        test_data[189] = 33'd257588625;
        test_addr[190] = 488;
        test_data[190] = 33'd2484186896;
        test_addr[191] = 958;
        test_data[191] = 33'd3257284543;
        test_addr[192] = 362;
        test_data[192] = 33'd4225808861;
        test_addr[193] = 855;
        test_data[193] = 33'd4260287046;
        test_addr[194] = 80;
        test_data[194] = 33'd818068638;
        test_addr[195] = 173;
        test_data[195] = 33'd1456155483;
        test_addr[196] = 584;
        test_data[196] = 33'd3681182924;
        test_addr[197] = 943;
        test_data[197] = 33'd7745382553;
        test_addr[198] = 114;
        test_data[198] = 33'd3614315923;
        test_addr[199] = 136;
        test_data[199] = 33'd3884710849;
        test_addr[200] = 66;
        test_data[200] = 33'd2051708468;
        test_addr[201] = 254;
        test_data[201] = 33'd4032840749;
        test_addr[202] = 416;
        test_data[202] = 33'd3819993292;
        test_addr[203] = 151;
        test_data[203] = 33'd199031358;
        test_addr[204] = 724;
        test_data[204] = 33'd8525596318;
        test_addr[205] = 235;
        test_data[205] = 33'd4802901797;
        test_addr[206] = 49;
        test_data[206] = 33'd751512591;
        test_addr[207] = 50;
        test_data[207] = 33'd5728089968;
        test_addr[208] = 975;
        test_data[208] = 33'd5981921165;
        test_addr[209] = 953;
        test_data[209] = 33'd5665203792;
        test_addr[210] = 657;
        test_data[210] = 33'd7815806751;
        test_addr[211] = 258;
        test_data[211] = 33'd7269271488;
        test_addr[212] = 313;
        test_data[212] = 33'd362309121;
        test_addr[213] = 5;
        test_data[213] = 33'd7058728075;
        test_addr[214] = 5;
        test_data[214] = 33'd2763760779;
        test_addr[215] = 444;
        test_data[215] = 33'd2124914818;
        test_addr[216] = 282;
        test_data[216] = 33'd8144760444;
        test_addr[217] = 813;
        test_data[217] = 33'd350957292;
        test_addr[218] = 278;
        test_data[218] = 33'd3400886719;
        test_addr[219] = 520;
        test_data[219] = 33'd3687095609;
        test_addr[220] = 660;
        test_data[220] = 33'd8341518676;
        test_addr[221] = 330;
        test_data[221] = 33'd2287195610;
        test_addr[222] = 1011;
        test_data[222] = 33'd6419460978;
        test_addr[223] = 984;
        test_data[223] = 33'd1155886029;
        test_addr[224] = 440;
        test_data[224] = 33'd5330839829;
        test_addr[225] = 334;
        test_data[225] = 33'd3431054307;
        test_addr[226] = 323;
        test_data[226] = 33'd5327415686;
        test_addr[227] = 797;
        test_data[227] = 33'd2090589244;
        test_addr[228] = 365;
        test_data[228] = 33'd369210451;
        test_addr[229] = 908;
        test_data[229] = 33'd1044409057;
        test_addr[230] = 665;
        test_data[230] = 33'd1128756264;
        test_addr[231] = 151;
        test_data[231] = 33'd7340079543;
        test_addr[232] = 273;
        test_data[232] = 33'd56693191;
        test_addr[233] = 175;
        test_data[233] = 33'd4957921855;
        test_addr[234] = 410;
        test_data[234] = 33'd3405405453;
        test_addr[235] = 88;
        test_data[235] = 33'd4094716213;
        test_addr[236] = 416;
        test_data[236] = 33'd3819993292;
        test_addr[237] = 288;
        test_data[237] = 33'd7961835817;
        test_addr[238] = 206;
        test_data[238] = 33'd380753888;
        test_addr[239] = 598;
        test_data[239] = 33'd3684002157;
        test_addr[240] = 700;
        test_data[240] = 33'd5054010116;
        test_addr[241] = 298;
        test_data[241] = 33'd1530159267;
        test_addr[242] = 747;
        test_data[242] = 33'd8562074142;
        test_addr[243] = 797;
        test_data[243] = 33'd2090589244;
        test_addr[244] = 320;
        test_data[244] = 33'd3248669603;
        test_addr[245] = 634;
        test_data[245] = 33'd2731773946;
        test_addr[246] = 239;
        test_data[246] = 33'd1377847727;
        test_addr[247] = 840;
        test_data[247] = 33'd8228101029;
        test_addr[248] = 347;
        test_data[248] = 33'd2552236765;
        test_addr[249] = 640;
        test_data[249] = 33'd7777171824;
        test_addr[250] = 952;
        test_data[250] = 33'd702855526;
        test_addr[251] = 239;
        test_data[251] = 33'd1377847727;
        test_addr[252] = 557;
        test_data[252] = 33'd7169721915;
        test_addr[253] = 676;
        test_data[253] = 33'd1174454579;
        test_addr[254] = 864;
        test_data[254] = 33'd1571587926;
        test_addr[255] = 20;
        test_data[255] = 33'd892044972;
        test_addr[256] = 59;
        test_data[256] = 33'd6219434332;
        test_addr[257] = 95;
        test_data[257] = 33'd3966602676;
        test_addr[258] = 244;
        test_data[258] = 33'd1306044194;
        test_addr[259] = 48;
        test_data[259] = 33'd8043244256;
        test_addr[260] = 196;
        test_data[260] = 33'd2957372585;
        test_addr[261] = 233;
        test_data[261] = 33'd1289878889;
        test_addr[262] = 94;
        test_data[262] = 33'd6786582673;
        test_addr[263] = 572;
        test_data[263] = 33'd2337695322;
        test_addr[264] = 404;
        test_data[264] = 33'd2626802031;
        test_addr[265] = 414;
        test_data[265] = 33'd402300966;
        test_addr[266] = 131;
        test_data[266] = 33'd813280569;
        test_addr[267] = 244;
        test_data[267] = 33'd4951927491;
        test_addr[268] = 111;
        test_data[268] = 33'd7757716555;
        test_addr[269] = 93;
        test_data[269] = 33'd263550839;
        test_addr[270] = 807;
        test_data[270] = 33'd4550572080;
        test_addr[271] = 775;
        test_data[271] = 33'd8559143006;
        test_addr[272] = 753;
        test_data[272] = 33'd7190779414;
        test_addr[273] = 532;
        test_data[273] = 33'd27322558;
        test_addr[274] = 804;
        test_data[274] = 33'd2469310094;
        test_addr[275] = 9;
        test_data[275] = 33'd5928931506;
        test_addr[276] = 164;
        test_data[276] = 33'd1777912528;
        test_addr[277] = 736;
        test_data[277] = 33'd6226581292;
        test_addr[278] = 222;
        test_data[278] = 33'd1146860549;
        test_addr[279] = 622;
        test_data[279] = 33'd7646389259;
        test_addr[280] = 416;
        test_data[280] = 33'd3819993292;
        test_addr[281] = 337;
        test_data[281] = 33'd1691010132;
        test_addr[282] = 626;
        test_data[282] = 33'd1808868451;
        test_addr[283] = 744;
        test_data[283] = 33'd7380109345;
        test_addr[284] = 135;
        test_data[284] = 33'd4364824501;
        test_addr[285] = 391;
        test_data[285] = 33'd2934085416;
        test_addr[286] = 924;
        test_data[286] = 33'd6059299042;
        test_addr[287] = 639;
        test_data[287] = 33'd382292317;
        test_addr[288] = 196;
        test_data[288] = 33'd5046070825;
        test_addr[289] = 71;
        test_data[289] = 33'd3950328245;
        test_addr[290] = 777;
        test_data[290] = 33'd485989889;
        test_addr[291] = 111;
        test_data[291] = 33'd3462749259;
        test_addr[292] = 604;
        test_data[292] = 33'd70723367;
        test_addr[293] = 513;
        test_data[293] = 33'd3717675145;
        test_addr[294] = 126;
        test_data[294] = 33'd2525024090;
        test_addr[295] = 55;
        test_data[295] = 33'd8584248253;
        test_addr[296] = 900;
        test_data[296] = 33'd8010696838;
        test_addr[297] = 576;
        test_data[297] = 33'd2373603425;
        test_addr[298] = 920;
        test_data[298] = 33'd3925196331;
        test_addr[299] = 702;
        test_data[299] = 33'd3866435097;
        test_addr[300] = 137;
        test_data[300] = 33'd1980778037;
        test_addr[301] = 602;
        test_data[301] = 33'd2312199791;
        test_addr[302] = 53;
        test_data[302] = 33'd4716342677;
        test_addr[303] = 673;
        test_data[303] = 33'd41814705;
        test_addr[304] = 848;
        test_data[304] = 33'd6281102252;
        test_addr[305] = 574;
        test_data[305] = 33'd2900017555;
        test_addr[306] = 800;
        test_data[306] = 33'd2470310901;
        test_addr[307] = 443;
        test_data[307] = 33'd8552951093;
        test_addr[308] = 924;
        test_data[308] = 33'd1764331746;
        test_addr[309] = 846;
        test_data[309] = 33'd2063463330;
        test_addr[310] = 790;
        test_data[310] = 33'd7263382786;
        test_addr[311] = 942;
        test_data[311] = 33'd4102784705;
        test_addr[312] = 588;
        test_data[312] = 33'd8336230681;
        test_addr[313] = 264;
        test_data[313] = 33'd687477629;
        test_addr[314] = 275;
        test_data[314] = 33'd8339129752;
        test_addr[315] = 948;
        test_data[315] = 33'd5011482461;
        test_addr[316] = 257;
        test_data[316] = 33'd894384987;
        test_addr[317] = 255;
        test_data[317] = 33'd6386041495;
        test_addr[318] = 715;
        test_data[318] = 33'd3660057142;
        test_addr[319] = 929;
        test_data[319] = 33'd2947338001;
        test_addr[320] = 110;
        test_data[320] = 33'd5211212181;
        test_addr[321] = 22;
        test_data[321] = 33'd9397193;
        test_addr[322] = 554;
        test_data[322] = 33'd302584709;
        test_addr[323] = 26;
        test_data[323] = 33'd6061194164;
        test_addr[324] = 638;
        test_data[324] = 33'd6991870293;
        test_addr[325] = 749;
        test_data[325] = 33'd5296534766;
        test_addr[326] = 43;
        test_data[326] = 33'd2636643983;
        test_addr[327] = 804;
        test_data[327] = 33'd2469310094;
        test_addr[328] = 873;
        test_data[328] = 33'd722926779;
        test_addr[329] = 908;
        test_data[329] = 33'd1044409057;
        test_addr[330] = 186;
        test_data[330] = 33'd4570927123;
        test_addr[331] = 841;
        test_data[331] = 33'd124879403;
        test_addr[332] = 938;
        test_data[332] = 33'd5854327783;
        test_addr[333] = 369;
        test_data[333] = 33'd1161521471;
        test_addr[334] = 367;
        test_data[334] = 33'd3620341239;
        test_addr[335] = 492;
        test_data[335] = 33'd2984910114;
        test_addr[336] = 350;
        test_data[336] = 33'd8271861287;
        test_addr[337] = 227;
        test_data[337] = 33'd905576619;
        test_addr[338] = 866;
        test_data[338] = 33'd3574629408;
        test_addr[339] = 216;
        test_data[339] = 33'd7339845595;
        test_addr[340] = 867;
        test_data[340] = 33'd18555133;
        test_addr[341] = 338;
        test_data[341] = 33'd3573453669;
        test_addr[342] = 960;
        test_data[342] = 33'd5405932872;
        test_addr[343] = 576;
        test_data[343] = 33'd6119941832;
        test_addr[344] = 274;
        test_data[344] = 33'd3318236443;
        test_addr[345] = 276;
        test_data[345] = 33'd2694496543;
        test_addr[346] = 363;
        test_data[346] = 33'd4960267679;
        test_addr[347] = 549;
        test_data[347] = 33'd8050293025;
        test_addr[348] = 466;
        test_data[348] = 33'd633115602;
        test_addr[349] = 1003;
        test_data[349] = 33'd5830313804;
        test_addr[350] = 33;
        test_data[350] = 33'd3931481952;
        test_addr[351] = 148;
        test_data[351] = 33'd3002299453;
        test_addr[352] = 301;
        test_data[352] = 33'd3075188539;
        test_addr[353] = 703;
        test_data[353] = 33'd4966731480;
        test_addr[354] = 571;
        test_data[354] = 33'd8144020506;
        test_addr[355] = 83;
        test_data[355] = 33'd681728304;
        test_addr[356] = 525;
        test_data[356] = 33'd426532196;
        test_addr[357] = 1003;
        test_data[357] = 33'd6415252152;
        test_addr[358] = 805;
        test_data[358] = 33'd692126376;
        test_addr[359] = 350;
        test_data[359] = 33'd3976893991;
        test_addr[360] = 997;
        test_data[360] = 33'd2903693877;
        test_addr[361] = 397;
        test_data[361] = 33'd2724761539;
        test_addr[362] = 881;
        test_data[362] = 33'd554101517;
        test_addr[363] = 560;
        test_data[363] = 33'd3890402307;
        test_addr[364] = 538;
        test_data[364] = 33'd1157057488;
        test_addr[365] = 679;
        test_data[365] = 33'd5768941855;
        test_addr[366] = 505;
        test_data[366] = 33'd5340133097;
        test_addr[367] = 210;
        test_data[367] = 33'd2782581352;
        test_addr[368] = 507;
        test_data[368] = 33'd3857079307;
        test_addr[369] = 652;
        test_data[369] = 33'd2524346705;
        test_addr[370] = 997;
        test_data[370] = 33'd5792842315;
        test_addr[371] = 890;
        test_data[371] = 33'd1689472630;
        test_addr[372] = 259;
        test_data[372] = 33'd3390847646;
        test_addr[373] = 303;
        test_data[373] = 33'd143048814;
        test_addr[374] = 883;
        test_data[374] = 33'd6090672700;
        test_addr[375] = 261;
        test_data[375] = 33'd629678269;
        test_addr[376] = 432;
        test_data[376] = 33'd926426471;
        test_addr[377] = 923;
        test_data[377] = 33'd6774514208;
        test_addr[378] = 602;
        test_data[378] = 33'd2312199791;
        test_addr[379] = 279;
        test_data[379] = 33'd6474833190;
        test_addr[380] = 82;
        test_data[380] = 33'd5568545962;
        test_addr[381] = 405;
        test_data[381] = 33'd6265027707;
        test_addr[382] = 55;
        test_data[382] = 33'd4289280957;
        test_addr[383] = 65;
        test_data[383] = 33'd993562414;
        test_addr[384] = 99;
        test_data[384] = 33'd2883454270;
        test_addr[385] = 66;
        test_data[385] = 33'd2051708468;
        test_addr[386] = 264;
        test_data[386] = 33'd687477629;
        test_addr[387] = 451;
        test_data[387] = 33'd317087304;
        test_addr[388] = 478;
        test_data[388] = 33'd627300334;
        test_addr[389] = 943;
        test_data[389] = 33'd8040433360;
        test_addr[390] = 339;
        test_data[390] = 33'd944678627;
        test_addr[391] = 39;
        test_data[391] = 33'd3097257097;
        test_addr[392] = 956;
        test_data[392] = 33'd6518506232;
        test_addr[393] = 430;
        test_data[393] = 33'd8207020564;
        test_addr[394] = 70;
        test_data[394] = 33'd1368704711;
        test_addr[395] = 209;
        test_data[395] = 33'd87559006;
        test_addr[396] = 722;
        test_data[396] = 33'd5940466549;
        test_addr[397] = 611;
        test_data[397] = 33'd2223272245;
        test_addr[398] = 789;
        test_data[398] = 33'd2899379877;
        test_addr[399] = 851;
        test_data[399] = 33'd550630034;
        test_addr[400] = 1003;
        test_data[400] = 33'd5578089764;
        test_addr[401] = 146;
        test_data[401] = 33'd2005652566;
        test_addr[402] = 207;
        test_data[402] = 33'd843754471;
        test_addr[403] = 834;
        test_data[403] = 33'd7477910575;
        test_addr[404] = 727;
        test_data[404] = 33'd2717525231;
        test_addr[405] = 734;
        test_data[405] = 33'd3464739256;
        test_addr[406] = 890;
        test_data[406] = 33'd6313394651;
        test_addr[407] = 263;
        test_data[407] = 33'd7577251992;
        test_addr[408] = 469;
        test_data[408] = 33'd7506568092;
        test_addr[409] = 1016;
        test_data[409] = 33'd6386386341;
        test_addr[410] = 941;
        test_data[410] = 33'd3244851306;
        test_addr[411] = 728;
        test_data[411] = 33'd128590783;
        test_addr[412] = 87;
        test_data[412] = 33'd2854372909;
        test_addr[413] = 931;
        test_data[413] = 33'd2803979244;
        test_addr[414] = 525;
        test_data[414] = 33'd426532196;
        test_addr[415] = 834;
        test_data[415] = 33'd3182943279;
        test_addr[416] = 421;
        test_data[416] = 33'd7394667507;
        test_addr[417] = 881;
        test_data[417] = 33'd554101517;
        test_addr[418] = 105;
        test_data[418] = 33'd3407001355;
        test_addr[419] = 749;
        test_data[419] = 33'd1001567470;
        test_addr[420] = 553;
        test_data[420] = 33'd4101269385;
        test_addr[421] = 294;
        test_data[421] = 33'd228860212;
        test_addr[422] = 780;
        test_data[422] = 33'd404411201;
        test_addr[423] = 707;
        test_data[423] = 33'd982366389;
        test_addr[424] = 337;
        test_data[424] = 33'd1691010132;
        test_addr[425] = 532;
        test_data[425] = 33'd7768145488;
        test_addr[426] = 898;
        test_data[426] = 33'd8359574126;
        test_addr[427] = 927;
        test_data[427] = 33'd1927721038;
        test_addr[428] = 108;
        test_data[428] = 33'd52659899;
        test_addr[429] = 789;
        test_data[429] = 33'd2899379877;
        test_addr[430] = 86;
        test_data[430] = 33'd7193033190;
        test_addr[431] = 812;
        test_data[431] = 33'd2625492882;
        test_addr[432] = 802;
        test_data[432] = 33'd6776085908;
        test_addr[433] = 918;
        test_data[433] = 33'd2681524291;
        test_addr[434] = 207;
        test_data[434] = 33'd843754471;
        test_addr[435] = 256;
        test_data[435] = 33'd5626177527;
        test_addr[436] = 647;
        test_data[436] = 33'd738418394;
        test_addr[437] = 1023;
        test_data[437] = 33'd4557021752;
        test_addr[438] = 315;
        test_data[438] = 33'd1263301752;
        test_addr[439] = 979;
        test_data[439] = 33'd1509757740;
        test_addr[440] = 247;
        test_data[440] = 33'd8303978359;
        test_addr[441] = 845;
        test_data[441] = 33'd6258713695;
        test_addr[442] = 920;
        test_data[442] = 33'd6130247968;
        test_addr[443] = 234;
        test_data[443] = 33'd8169106890;
        test_addr[444] = 832;
        test_data[444] = 33'd351971474;
        test_addr[445] = 10;
        test_data[445] = 33'd4085122833;
        test_addr[446] = 28;
        test_data[446] = 33'd1087055728;
        test_addr[447] = 788;
        test_data[447] = 33'd3121816568;
        test_addr[448] = 517;
        test_data[448] = 33'd385111081;
        test_addr[449] = 167;
        test_data[449] = 33'd188544578;
        test_addr[450] = 46;
        test_data[450] = 33'd1936612333;
        test_addr[451] = 854;
        test_data[451] = 33'd2260897852;
        test_addr[452] = 18;
        test_data[452] = 33'd7665762087;
        test_addr[453] = 0;
        test_data[453] = 33'd3214325899;
        test_addr[454] = 390;
        test_data[454] = 33'd909123417;
        test_addr[455] = 984;
        test_data[455] = 33'd1155886029;
        test_addr[456] = 965;
        test_data[456] = 33'd7861830793;
        test_addr[457] = 921;
        test_data[457] = 33'd680034433;
        test_addr[458] = 507;
        test_data[458] = 33'd3857079307;
        test_addr[459] = 532;
        test_data[459] = 33'd3473178192;
        test_addr[460] = 870;
        test_data[460] = 33'd4461659300;
        test_addr[461] = 318;
        test_data[461] = 33'd5513831788;
        test_addr[462] = 636;
        test_data[462] = 33'd3726205383;
        test_addr[463] = 178;
        test_data[463] = 33'd3283596447;
        test_addr[464] = 77;
        test_data[464] = 33'd1279103495;
        test_addr[465] = 82;
        test_data[465] = 33'd7403099325;
        test_addr[466] = 568;
        test_data[466] = 33'd2796273124;
        test_addr[467] = 674;
        test_data[467] = 33'd2656360569;
        test_addr[468] = 160;
        test_data[468] = 33'd1681817037;
        test_addr[469] = 139;
        test_data[469] = 33'd8476938710;
        test_addr[470] = 39;
        test_data[470] = 33'd3097257097;
        test_addr[471] = 960;
        test_data[471] = 33'd1110965576;
        test_addr[472] = 635;
        test_data[472] = 33'd604312534;
        test_addr[473] = 236;
        test_data[473] = 33'd983334167;
        test_addr[474] = 154;
        test_data[474] = 33'd1881539630;
        test_addr[475] = 844;
        test_data[475] = 33'd1272998109;
        test_addr[476] = 929;
        test_data[476] = 33'd2947338001;
        test_addr[477] = 125;
        test_data[477] = 33'd2709632180;
        test_addr[478] = 328;
        test_data[478] = 33'd952282828;
        test_addr[479] = 259;
        test_data[479] = 33'd3390847646;
        test_addr[480] = 594;
        test_data[480] = 33'd3790697293;
        test_addr[481] = 773;
        test_data[481] = 33'd2884864817;
        test_addr[482] = 876;
        test_data[482] = 33'd7217237352;
        test_addr[483] = 585;
        test_data[483] = 33'd3586969900;
        test_addr[484] = 466;
        test_data[484] = 33'd633115602;
        test_addr[485] = 750;
        test_data[485] = 33'd4675191772;
        test_addr[486] = 389;
        test_data[486] = 33'd2549642068;
        test_addr[487] = 1005;
        test_data[487] = 33'd1098300837;
        test_addr[488] = 553;
        test_data[488] = 33'd4101269385;
        test_addr[489] = 547;
        test_data[489] = 33'd7395375881;
        test_addr[490] = 937;
        test_data[490] = 33'd3186542920;
        test_addr[491] = 633;
        test_data[491] = 33'd6081308139;
        test_addr[492] = 708;
        test_data[492] = 33'd7658518223;
        test_addr[493] = 545;
        test_data[493] = 33'd3465705991;
        test_addr[494] = 104;
        test_data[494] = 33'd3714367826;
        test_addr[495] = 409;
        test_data[495] = 33'd5608659419;
        test_addr[496] = 502;
        test_data[496] = 33'd6172771661;
        test_addr[497] = 648;
        test_data[497] = 33'd6320829636;
        test_addr[498] = 520;
        test_data[498] = 33'd8436810523;
        test_addr[499] = 640;
        test_data[499] = 33'd3482204528;
        test_addr[500] = 248;
        test_data[500] = 33'd810408981;
        test_addr[501] = 751;
        test_data[501] = 33'd7018041834;
        test_addr[502] = 29;
        test_data[502] = 33'd4426040515;
        test_addr[503] = 66;
        test_data[503] = 33'd2051708468;
        test_addr[504] = 10;
        test_data[504] = 33'd4085122833;
        test_addr[505] = 208;
        test_data[505] = 33'd5834224912;
        test_addr[506] = 397;
        test_data[506] = 33'd6786474336;
        test_addr[507] = 582;
        test_data[507] = 33'd7063246473;
        test_addr[508] = 4;
        test_data[508] = 33'd5612750778;
        test_addr[509] = 534;
        test_data[509] = 33'd5013108132;
        test_addr[510] = 592;
        test_data[510] = 33'd3006473031;
        test_addr[511] = 877;
        test_data[511] = 33'd5134426982;
        test_addr[512] = 496;
        test_data[512] = 33'd1048502686;
        test_addr[513] = 673;
        test_data[513] = 33'd41814705;
        test_addr[514] = 1021;
        test_data[514] = 33'd707276233;
        test_addr[515] = 655;
        test_data[515] = 33'd2678884701;
        test_addr[516] = 836;
        test_data[516] = 33'd1052769268;
        test_addr[517] = 126;
        test_data[517] = 33'd2525024090;
        test_addr[518] = 511;
        test_data[518] = 33'd308446067;
        test_addr[519] = 992;
        test_data[519] = 33'd7578883622;
        test_addr[520] = 467;
        test_data[520] = 33'd3833383596;
        test_addr[521] = 497;
        test_data[521] = 33'd2590240532;
        test_addr[522] = 237;
        test_data[522] = 33'd2066899154;
        test_addr[523] = 114;
        test_data[523] = 33'd3614315923;
        test_addr[524] = 206;
        test_data[524] = 33'd380753888;
        test_addr[525] = 0;
        test_data[525] = 33'd3214325899;
        test_addr[526] = 164;
        test_data[526] = 33'd1777912528;
        test_addr[527] = 1021;
        test_data[527] = 33'd7765783293;
        test_addr[528] = 161;
        test_data[528] = 33'd7936775649;
        test_addr[529] = 33;
        test_data[529] = 33'd7215764017;
        test_addr[530] = 7;
        test_data[530] = 33'd881802803;
        test_addr[531] = 506;
        test_data[531] = 33'd644403250;
        test_addr[532] = 242;
        test_data[532] = 33'd6277782442;
        test_addr[533] = 735;
        test_data[533] = 33'd8482548222;
        test_addr[534] = 681;
        test_data[534] = 33'd1893449825;
        test_addr[535] = 830;
        test_data[535] = 33'd5864876069;
        test_addr[536] = 930;
        test_data[536] = 33'd6302525038;
        test_addr[537] = 922;
        test_data[537] = 33'd715587172;
        test_addr[538] = 315;
        test_data[538] = 33'd1263301752;
        test_addr[539] = 103;
        test_data[539] = 33'd2627891325;
        test_addr[540] = 459;
        test_data[540] = 33'd8545729866;
        test_addr[541] = 274;
        test_data[541] = 33'd3318236443;
        test_addr[542] = 509;
        test_data[542] = 33'd1404134308;
        test_addr[543] = 647;
        test_data[543] = 33'd4301913415;
        test_addr[544] = 446;
        test_data[544] = 33'd3099163608;
        test_addr[545] = 59;
        test_data[545] = 33'd1924467036;
        test_addr[546] = 556;
        test_data[546] = 33'd6325765236;
        test_addr[547] = 974;
        test_data[547] = 33'd2073535736;
        test_addr[548] = 176;
        test_data[548] = 33'd2275341057;
        test_addr[549] = 467;
        test_data[549] = 33'd7223830261;
        test_addr[550] = 275;
        test_data[550] = 33'd4044162456;
        test_addr[551] = 432;
        test_data[551] = 33'd5563554304;
        test_addr[552] = 168;
        test_data[552] = 33'd4914390344;
        test_addr[553] = 97;
        test_data[553] = 33'd2839264634;
        test_addr[554] = 991;
        test_data[554] = 33'd3554038044;
        test_addr[555] = 286;
        test_data[555] = 33'd2360048588;
        test_addr[556] = 965;
        test_data[556] = 33'd3566863497;
        test_addr[557] = 267;
        test_data[557] = 33'd3627326475;
        test_addr[558] = 127;
        test_data[558] = 33'd6026400207;
        test_addr[559] = 138;
        test_data[559] = 33'd2910298998;
        test_addr[560] = 427;
        test_data[560] = 33'd3998550133;
        test_addr[561] = 880;
        test_data[561] = 33'd1923216062;
        test_addr[562] = 370;
        test_data[562] = 33'd5834892018;
        test_addr[563] = 873;
        test_data[563] = 33'd722926779;
        test_addr[564] = 59;
        test_data[564] = 33'd1924467036;
        test_addr[565] = 370;
        test_data[565] = 33'd1539924722;
        test_addr[566] = 202;
        test_data[566] = 33'd7055529581;
        test_addr[567] = 814;
        test_data[567] = 33'd662516995;
        test_addr[568] = 107;
        test_data[568] = 33'd4243198286;
        test_addr[569] = 192;
        test_data[569] = 33'd2694434016;
        test_addr[570] = 119;
        test_data[570] = 33'd1052542082;
        test_addr[571] = 921;
        test_data[571] = 33'd8297010819;
        test_addr[572] = 746;
        test_data[572] = 33'd2332255621;
        test_addr[573] = 101;
        test_data[573] = 33'd5126825292;
        test_addr[574] = 776;
        test_data[574] = 33'd769284591;
        test_addr[575] = 458;
        test_data[575] = 33'd3114864730;
        test_addr[576] = 582;
        test_data[576] = 33'd6222658799;
        test_addr[577] = 215;
        test_data[577] = 33'd7466796527;
        test_addr[578] = 277;
        test_data[578] = 33'd7094759426;
        test_addr[579] = 87;
        test_data[579] = 33'd2854372909;
        test_addr[580] = 356;
        test_data[580] = 33'd2587005368;
        test_addr[581] = 682;
        test_data[581] = 33'd4596873333;
        test_addr[582] = 846;
        test_data[582] = 33'd2063463330;
        test_addr[583] = 937;
        test_data[583] = 33'd3186542920;
        test_addr[584] = 177;
        test_data[584] = 33'd2198187797;
        test_addr[585] = 710;
        test_data[585] = 33'd4248041353;
        test_addr[586] = 673;
        test_data[586] = 33'd41814705;
        test_addr[587] = 196;
        test_data[587] = 33'd751103529;
        test_addr[588] = 10;
        test_data[588] = 33'd7889776412;
        test_addr[589] = 429;
        test_data[589] = 33'd3992289899;
        test_addr[590] = 496;
        test_data[590] = 33'd4777640912;
        test_addr[591] = 706;
        test_data[591] = 33'd5080209594;
        test_addr[592] = 507;
        test_data[592] = 33'd3857079307;
        test_addr[593] = 391;
        test_data[593] = 33'd2934085416;
        test_addr[594] = 974;
        test_data[594] = 33'd2073535736;
        test_addr[595] = 17;
        test_data[595] = 33'd2023586953;
        test_addr[596] = 908;
        test_data[596] = 33'd5429599875;
        test_addr[597] = 35;
        test_data[597] = 33'd1427007413;
        test_addr[598] = 734;
        test_data[598] = 33'd3464739256;
        test_addr[599] = 190;
        test_data[599] = 33'd2487141371;
        test_addr[600] = 608;
        test_data[600] = 33'd3381739994;
        test_addr[601] = 513;
        test_data[601] = 33'd3717675145;
        test_addr[602] = 194;
        test_data[602] = 33'd2912051046;
        test_addr[603] = 315;
        test_data[603] = 33'd1263301752;
        test_addr[604] = 811;
        test_data[604] = 33'd712960676;
        test_addr[605] = 499;
        test_data[605] = 33'd4266444285;
        test_addr[606] = 608;
        test_data[606] = 33'd3381739994;
        test_addr[607] = 946;
        test_data[607] = 33'd6084424548;
        test_addr[608] = 519;
        test_data[608] = 33'd1283402259;
        test_addr[609] = 719;
        test_data[609] = 33'd8075731471;
        test_addr[610] = 852;
        test_data[610] = 33'd6891579326;
        test_addr[611] = 706;
        test_data[611] = 33'd785242298;
        test_addr[612] = 920;
        test_data[612] = 33'd1835280672;
        test_addr[613] = 239;
        test_data[613] = 33'd1377847727;
        test_addr[614] = 209;
        test_data[614] = 33'd6823727363;
        test_addr[615] = 330;
        test_data[615] = 33'd2287195610;
        test_addr[616] = 191;
        test_data[616] = 33'd1599404350;
        test_addr[617] = 960;
        test_data[617] = 33'd5790857860;
        test_addr[618] = 960;
        test_data[618] = 33'd1495890564;
        test_addr[619] = 815;
        test_data[619] = 33'd1640602374;
        test_addr[620] = 208;
        test_data[620] = 33'd1539257616;
        test_addr[621] = 672;
        test_data[621] = 33'd3252626599;
        test_addr[622] = 972;
        test_data[622] = 33'd7872786849;
        test_addr[623] = 390;
        test_data[623] = 33'd909123417;
        test_addr[624] = 536;
        test_data[624] = 33'd2903832397;
        test_addr[625] = 731;
        test_data[625] = 33'd1134545885;
        test_addr[626] = 95;
        test_data[626] = 33'd3966602676;
        test_addr[627] = 675;
        test_data[627] = 33'd140747614;
        test_addr[628] = 787;
        test_data[628] = 33'd1935616810;
        test_addr[629] = 403;
        test_data[629] = 33'd6646913738;
        test_addr[630] = 508;
        test_data[630] = 33'd2569124247;
        test_addr[631] = 237;
        test_data[631] = 33'd2066899154;
        test_addr[632] = 1021;
        test_data[632] = 33'd3470815997;
        test_addr[633] = 7;
        test_data[633] = 33'd881802803;
        test_addr[634] = 95;
        test_data[634] = 33'd3966602676;
        test_addr[635] = 772;
        test_data[635] = 33'd3678900751;
        test_addr[636] = 372;
        test_data[636] = 33'd3706783982;
        test_addr[637] = 82;
        test_data[637] = 33'd5475737146;
        test_addr[638] = 580;
        test_data[638] = 33'd436662051;
        test_addr[639] = 225;
        test_data[639] = 33'd541535233;
        test_addr[640] = 489;
        test_data[640] = 33'd5537091895;
        test_addr[641] = 354;
        test_data[641] = 33'd2820300650;
        test_addr[642] = 705;
        test_data[642] = 33'd1506519041;
        test_addr[643] = 343;
        test_data[643] = 33'd2472167151;
        test_addr[644] = 531;
        test_data[644] = 33'd3479564107;
        test_addr[645] = 841;
        test_data[645] = 33'd124879403;
        test_addr[646] = 740;
        test_data[646] = 33'd2129383015;
        test_addr[647] = 271;
        test_data[647] = 33'd2718986291;
        test_addr[648] = 770;
        test_data[648] = 33'd5245554392;
        test_addr[649] = 197;
        test_data[649] = 33'd6688331653;
        test_addr[650] = 463;
        test_data[650] = 33'd1603013143;
        test_addr[651] = 1017;
        test_data[651] = 33'd7339940083;
        test_addr[652] = 378;
        test_data[652] = 33'd2059550719;
        test_addr[653] = 878;
        test_data[653] = 33'd1973087823;
        test_addr[654] = 681;
        test_data[654] = 33'd1893449825;
        test_addr[655] = 537;
        test_data[655] = 33'd810473933;
        test_addr[656] = 206;
        test_data[656] = 33'd380753888;
        test_addr[657] = 534;
        test_data[657] = 33'd6759855210;
        test_addr[658] = 174;
        test_data[658] = 33'd7899067612;
        test_addr[659] = 12;
        test_data[659] = 33'd4028186270;
        test_addr[660] = 878;
        test_data[660] = 33'd4769728491;
        test_addr[661] = 100;
        test_data[661] = 33'd3239304748;
        test_addr[662] = 489;
        test_data[662] = 33'd1242124599;
        test_addr[663] = 986;
        test_data[663] = 33'd6376562981;
        test_addr[664] = 450;
        test_data[664] = 33'd2461350224;
        test_addr[665] = 735;
        test_data[665] = 33'd4187580926;
        test_addr[666] = 639;
        test_data[666] = 33'd8492686316;
        test_addr[667] = 257;
        test_data[667] = 33'd894384987;
        test_addr[668] = 793;
        test_data[668] = 33'd1650429696;
        test_addr[669] = 910;
        test_data[669] = 33'd4293745703;
        test_addr[670] = 201;
        test_data[670] = 33'd29735866;
        test_addr[671] = 422;
        test_data[671] = 33'd4144807526;
        test_addr[672] = 414;
        test_data[672] = 33'd402300966;
        test_addr[673] = 458;
        test_data[673] = 33'd3114864730;
        test_addr[674] = 333;
        test_data[674] = 33'd509475252;
        test_addr[675] = 505;
        test_data[675] = 33'd1045165801;
        test_addr[676] = 67;
        test_data[676] = 33'd3639768664;
        test_addr[677] = 554;
        test_data[677] = 33'd302584709;
        test_addr[678] = 328;
        test_data[678] = 33'd952282828;
        test_addr[679] = 773;
        test_data[679] = 33'd5437894622;
        test_addr[680] = 497;
        test_data[680] = 33'd5279502434;
        test_addr[681] = 397;
        test_data[681] = 33'd2491507040;
        test_addr[682] = 803;
        test_data[682] = 33'd1913165819;
        test_addr[683] = 562;
        test_data[683] = 33'd8403921312;
        test_addr[684] = 555;
        test_data[684] = 33'd920282072;
        test_addr[685] = 715;
        test_data[685] = 33'd3660057142;
        test_addr[686] = 831;
        test_data[686] = 33'd992727670;
        test_addr[687] = 627;
        test_data[687] = 33'd1310702174;
        test_addr[688] = 590;
        test_data[688] = 33'd6002574066;
        test_addr[689] = 729;
        test_data[689] = 33'd1035742076;
        test_addr[690] = 592;
        test_data[690] = 33'd5233760978;
        test_addr[691] = 166;
        test_data[691] = 33'd5512843665;
        test_addr[692] = 658;
        test_data[692] = 33'd1232299630;
        test_addr[693] = 20;
        test_data[693] = 33'd892044972;
        test_addr[694] = 107;
        test_data[694] = 33'd4243198286;
        test_addr[695] = 43;
        test_data[695] = 33'd2636643983;
        test_addr[696] = 10;
        test_data[696] = 33'd3594809116;
        test_addr[697] = 268;
        test_data[697] = 33'd59643427;
        test_addr[698] = 63;
        test_data[698] = 33'd100769450;
        test_addr[699] = 647;
        test_data[699] = 33'd6946119;
        test_addr[700] = 707;
        test_data[700] = 33'd6746348287;
        test_addr[701] = 489;
        test_data[701] = 33'd1242124599;
        test_addr[702] = 421;
        test_data[702] = 33'd8438354433;
        test_addr[703] = 146;
        test_data[703] = 33'd7734992814;
        test_addr[704] = 554;
        test_data[704] = 33'd6502151062;
        test_addr[705] = 847;
        test_data[705] = 33'd196428976;
        test_addr[706] = 499;
        test_data[706] = 33'd4266444285;
        test_addr[707] = 906;
        test_data[707] = 33'd5827587084;
        test_addr[708] = 57;
        test_data[708] = 33'd2855835886;
        test_addr[709] = 939;
        test_data[709] = 33'd536731119;
        test_addr[710] = 42;
        test_data[710] = 33'd3652372969;
        test_addr[711] = 58;
        test_data[711] = 33'd8481234607;
        test_addr[712] = 812;
        test_data[712] = 33'd5406055263;
        test_addr[713] = 486;
        test_data[713] = 33'd2789818792;
        test_addr[714] = 239;
        test_data[714] = 33'd1377847727;
        test_addr[715] = 31;
        test_data[715] = 33'd1855015640;
        test_addr[716] = 793;
        test_data[716] = 33'd1650429696;
        test_addr[717] = 871;
        test_data[717] = 33'd3173545540;
        test_addr[718] = 920;
        test_data[718] = 33'd1835280672;
        test_addr[719] = 725;
        test_data[719] = 33'd5642364353;
        test_addr[720] = 175;
        test_data[720] = 33'd662954559;
        test_addr[721] = 959;
        test_data[721] = 33'd3913949685;
        test_addr[722] = 238;
        test_data[722] = 33'd5515050210;
        test_addr[723] = 920;
        test_data[723] = 33'd1835280672;
        test_addr[724] = 228;
        test_data[724] = 33'd3498918036;
        test_addr[725] = 6;
        test_data[725] = 33'd1280683540;
        test_addr[726] = 157;
        test_data[726] = 33'd7779355172;
        test_addr[727] = 1023;
        test_data[727] = 33'd262054456;
        test_addr[728] = 832;
        test_data[728] = 33'd351971474;
        test_addr[729] = 639;
        test_data[729] = 33'd4197719020;
        test_addr[730] = 312;
        test_data[730] = 33'd1985873362;
        test_addr[731] = 265;
        test_data[731] = 33'd8097730453;
        test_addr[732] = 984;
        test_data[732] = 33'd5719746040;
        test_addr[733] = 827;
        test_data[733] = 33'd4136395276;
        test_addr[734] = 611;
        test_data[734] = 33'd5098653155;
        test_addr[735] = 558;
        test_data[735] = 33'd3650811963;
        test_addr[736] = 841;
        test_data[736] = 33'd124879403;
        test_addr[737] = 871;
        test_data[737] = 33'd8195342212;
        test_addr[738] = 122;
        test_data[738] = 33'd1522076612;
        test_addr[739] = 119;
        test_data[739] = 33'd7058201621;
        test_addr[740] = 250;
        test_data[740] = 33'd673588786;
        test_addr[741] = 368;
        test_data[741] = 33'd3346930613;
        test_addr[742] = 835;
        test_data[742] = 33'd3461985819;
        test_addr[743] = 175;
        test_data[743] = 33'd662954559;
        test_addr[744] = 277;
        test_data[744] = 33'd2799792130;
        test_addr[745] = 534;
        test_data[745] = 33'd2464887914;
        test_addr[746] = 874;
        test_data[746] = 33'd2931664417;
        test_addr[747] = 283;
        test_data[747] = 33'd4875977297;
        test_addr[748] = 431;
        test_data[748] = 33'd3304810659;
        test_addr[749] = 469;
        test_data[749] = 33'd3211600796;
        test_addr[750] = 818;
        test_data[750] = 33'd8167456569;
        test_addr[751] = 0;
        test_data[751] = 33'd3214325899;
        test_addr[752] = 863;
        test_data[752] = 33'd1325550564;
        test_addr[753] = 688;
        test_data[753] = 33'd4133517367;
        test_addr[754] = 179;
        test_data[754] = 33'd3433493149;
        test_addr[755] = 195;
        test_data[755] = 33'd5309705343;
        test_addr[756] = 415;
        test_data[756] = 33'd330435490;
        test_addr[757] = 980;
        test_data[757] = 33'd2435006134;
        test_addr[758] = 310;
        test_data[758] = 33'd3692301779;
        test_addr[759] = 379;
        test_data[759] = 33'd7249400730;
        test_addr[760] = 77;
        test_data[760] = 33'd4518573081;
        test_addr[761] = 39;
        test_data[761] = 33'd3097257097;
        test_addr[762] = 103;
        test_data[762] = 33'd2627891325;
        test_addr[763] = 967;
        test_data[763] = 33'd3880369406;
        test_addr[764] = 240;
        test_data[764] = 33'd3107113144;
        test_addr[765] = 66;
        test_data[765] = 33'd2051708468;
        test_addr[766] = 21;
        test_data[766] = 33'd6009152391;
        test_addr[767] = 388;
        test_data[767] = 33'd5095957581;
        test_addr[768] = 574;
        test_data[768] = 33'd6624050010;
        test_addr[769] = 378;
        test_data[769] = 33'd7424710498;
        test_addr[770] = 998;
        test_data[770] = 33'd8192191660;
        test_addr[771] = 184;
        test_data[771] = 33'd3840564828;
        test_addr[772] = 213;
        test_data[772] = 33'd2155161093;
        test_addr[773] = 577;
        test_data[773] = 33'd831046106;
        test_addr[774] = 499;
        test_data[774] = 33'd6413577625;
        test_addr[775] = 215;
        test_data[775] = 33'd7698190530;
        test_addr[776] = 417;
        test_data[776] = 33'd2268883569;
        test_addr[777] = 638;
        test_data[777] = 33'd6450550222;
        test_addr[778] = 986;
        test_data[778] = 33'd2081595685;
        test_addr[779] = 29;
        test_data[779] = 33'd131073219;
        test_addr[780] = 524;
        test_data[780] = 33'd1899487675;
        test_addr[781] = 787;
        test_data[781] = 33'd1935616810;
        test_addr[782] = 178;
        test_data[782] = 33'd3283596447;
        test_addr[783] = 871;
        test_data[783] = 33'd3900374916;
        test_addr[784] = 518;
        test_data[784] = 33'd856602084;
        test_addr[785] = 533;
        test_data[785] = 33'd8103984541;
        test_addr[786] = 404;
        test_data[786] = 33'd2626802031;
        test_addr[787] = 33;
        test_data[787] = 33'd2920796721;
        test_addr[788] = 255;
        test_data[788] = 33'd7660762152;
        test_addr[789] = 584;
        test_data[789] = 33'd3681182924;
        test_addr[790] = 828;
        test_data[790] = 33'd4550461102;
        test_addr[791] = 507;
        test_data[791] = 33'd3857079307;
        test_addr[792] = 202;
        test_data[792] = 33'd2760562285;
        test_addr[793] = 699;
        test_data[793] = 33'd716758767;
        test_addr[794] = 543;
        test_data[794] = 33'd7664293657;
        test_addr[795] = 393;
        test_data[795] = 33'd7530434122;
        test_addr[796] = 561;
        test_data[796] = 33'd5645491918;
        test_addr[797] = 738;
        test_data[797] = 33'd1085936134;
        test_addr[798] = 640;
        test_data[798] = 33'd3482204528;
        test_addr[799] = 703;
        test_data[799] = 33'd671764184;
        test_addr[800] = 833;
        test_data[800] = 33'd5188269229;
        test_addr[801] = 720;
        test_data[801] = 33'd2954885626;
        test_addr[802] = 450;
        test_data[802] = 33'd2461350224;
        test_addr[803] = 1004;
        test_data[803] = 33'd7922528203;
        test_addr[804] = 815;
        test_data[804] = 33'd1640602374;
        test_addr[805] = 1013;
        test_data[805] = 33'd519919884;
        test_addr[806] = 837;
        test_data[806] = 33'd7315427255;
        test_addr[807] = 565;
        test_data[807] = 33'd2843637762;
        test_addr[808] = 652;
        test_data[808] = 33'd2524346705;
        test_addr[809] = 963;
        test_data[809] = 33'd2423315520;
        test_addr[810] = 460;
        test_data[810] = 33'd5841282911;
        test_addr[811] = 521;
        test_data[811] = 33'd3462858656;
        test_addr[812] = 803;
        test_data[812] = 33'd1913165819;
        test_addr[813] = 287;
        test_data[813] = 33'd3189797644;
        test_addr[814] = 525;
        test_data[814] = 33'd8127952950;
        test_addr[815] = 924;
        test_data[815] = 33'd1764331746;
        test_addr[816] = 396;
        test_data[816] = 33'd7070731353;
        test_addr[817] = 752;
        test_data[817] = 33'd811875741;
        test_addr[818] = 586;
        test_data[818] = 33'd3378604480;
        test_addr[819] = 475;
        test_data[819] = 33'd2883836476;
        test_addr[820] = 849;
        test_data[820] = 33'd5616674377;
        test_addr[821] = 165;
        test_data[821] = 33'd106644142;
        test_addr[822] = 685;
        test_data[822] = 33'd4026500536;
        test_addr[823] = 553;
        test_data[823] = 33'd8083390038;
        test_addr[824] = 964;
        test_data[824] = 33'd1077138145;
        test_addr[825] = 361;
        test_data[825] = 33'd7739686333;
        test_addr[826] = 795;
        test_data[826] = 33'd5495737865;
        test_addr[827] = 582;
        test_data[827] = 33'd1927691503;
        test_addr[828] = 1004;
        test_data[828] = 33'd3627560907;
        test_addr[829] = 200;
        test_data[829] = 33'd4007449550;
        test_addr[830] = 662;
        test_data[830] = 33'd6478746656;
        test_addr[831] = 61;
        test_data[831] = 33'd3243858099;
        test_addr[832] = 81;
        test_data[832] = 33'd3391775223;
        test_addr[833] = 944;
        test_data[833] = 33'd5057634370;
        test_addr[834] = 679;
        test_data[834] = 33'd1473974559;
        test_addr[835] = 554;
        test_data[835] = 33'd2207183766;
        test_addr[836] = 711;
        test_data[836] = 33'd2297538283;
        test_addr[837] = 946;
        test_data[837] = 33'd1789457252;
        test_addr[838] = 671;
        test_data[838] = 33'd565008109;
        test_addr[839] = 695;
        test_data[839] = 33'd2186911345;
        test_addr[840] = 492;
        test_data[840] = 33'd2984910114;
        test_addr[841] = 520;
        test_data[841] = 33'd8207563406;
        test_addr[842] = 4;
        test_data[842] = 33'd1317783482;
        test_addr[843] = 339;
        test_data[843] = 33'd944678627;
        test_addr[844] = 324;
        test_data[844] = 33'd330852185;
        test_addr[845] = 137;
        test_data[845] = 33'd5510502815;
        test_addr[846] = 516;
        test_data[846] = 33'd1259652408;
        test_addr[847] = 167;
        test_data[847] = 33'd188544578;
        test_addr[848] = 153;
        test_data[848] = 33'd632865373;
        test_addr[849] = 163;
        test_data[849] = 33'd1640167561;
        test_addr[850] = 139;
        test_data[850] = 33'd4181971414;
        test_addr[851] = 325;
        test_data[851] = 33'd539824620;
        test_addr[852] = 527;
        test_data[852] = 33'd1169423377;
        test_addr[853] = 41;
        test_data[853] = 33'd190445736;
        test_addr[854] = 650;
        test_data[854] = 33'd2885272839;
        test_addr[855] = 531;
        test_data[855] = 33'd3479564107;
        test_addr[856] = 681;
        test_data[856] = 33'd1893449825;
        test_addr[857] = 874;
        test_data[857] = 33'd2931664417;
        test_addr[858] = 820;
        test_data[858] = 33'd4175331955;
        test_addr[859] = 368;
        test_data[859] = 33'd3346930613;
        test_addr[860] = 132;
        test_data[860] = 33'd3529417599;
        test_addr[861] = 300;
        test_data[861] = 33'd5694534096;
        test_addr[862] = 273;
        test_data[862] = 33'd56693191;
        test_addr[863] = 60;
        test_data[863] = 33'd7190672408;
        test_addr[864] = 150;
        test_data[864] = 33'd1321807965;
        test_addr[865] = 777;
        test_data[865] = 33'd485989889;
        test_addr[866] = 557;
        test_data[866] = 33'd2874754619;
        test_addr[867] = 912;
        test_data[867] = 33'd1978461553;
        test_addr[868] = 720;
        test_data[868] = 33'd5008811917;
        test_addr[869] = 338;
        test_data[869] = 33'd7537550112;
        test_addr[870] = 602;
        test_data[870] = 33'd2312199791;
        test_addr[871] = 471;
        test_data[871] = 33'd1336088425;
        test_addr[872] = 602;
        test_data[872] = 33'd5341364892;
        test_addr[873] = 791;
        test_data[873] = 33'd2834578210;
        test_addr[874] = 350;
        test_data[874] = 33'd3976893991;
        test_addr[875] = 465;
        test_data[875] = 33'd5191787608;
        test_addr[876] = 82;
        test_data[876] = 33'd1180769850;
        test_addr[877] = 777;
        test_data[877] = 33'd485989889;
        test_addr[878] = 49;
        test_data[878] = 33'd751512591;
        test_addr[879] = 348;
        test_data[879] = 33'd6278973688;
        test_addr[880] = 794;
        test_data[880] = 33'd5753179239;
        test_addr[881] = 251;
        test_data[881] = 33'd1773791810;
        test_addr[882] = 775;
        test_data[882] = 33'd4264175710;
        test_addr[883] = 438;
        test_data[883] = 33'd2860390341;
        test_addr[884] = 834;
        test_data[884] = 33'd6081430408;
        test_addr[885] = 463;
        test_data[885] = 33'd1603013143;
        test_addr[886] = 971;
        test_data[886] = 33'd634864571;
        test_addr[887] = 858;
        test_data[887] = 33'd7549554987;
        test_addr[888] = 601;
        test_data[888] = 33'd2919076942;
        test_addr[889] = 899;
        test_data[889] = 33'd3868985293;
        test_addr[890] = 525;
        test_data[890] = 33'd6923950108;
        test_addr[891] = 451;
        test_data[891] = 33'd317087304;
        test_addr[892] = 27;
        test_data[892] = 33'd3441740048;
        test_addr[893] = 292;
        test_data[893] = 33'd2039041372;
        test_addr[894] = 650;
        test_data[894] = 33'd2885272839;
        test_addr[895] = 986;
        test_data[895] = 33'd2081595685;
        test_addr[896] = 599;
        test_data[896] = 33'd7782954771;
        test_addr[897] = 216;
        test_data[897] = 33'd3044878299;
        test_addr[898] = 996;
        test_data[898] = 33'd8070136648;
        test_addr[899] = 758;
        test_data[899] = 33'd879054465;
        test_addr[900] = 717;
        test_data[900] = 33'd2912310291;
        test_addr[901] = 245;
        test_data[901] = 33'd2052459312;
        test_addr[902] = 376;
        test_data[902] = 33'd3017136644;
        test_addr[903] = 229;
        test_data[903] = 33'd5215593745;
        test_addr[904] = 717;
        test_data[904] = 33'd7121231621;
        test_addr[905] = 742;
        test_data[905] = 33'd2915364435;
        test_addr[906] = 405;
        test_data[906] = 33'd4811076934;
        test_addr[907] = 536;
        test_data[907] = 33'd5972784173;
        test_addr[908] = 1016;
        test_data[908] = 33'd2091419045;
        test_addr[909] = 335;
        test_data[909] = 33'd7856294698;
        test_addr[910] = 164;
        test_data[910] = 33'd1777912528;
        test_addr[911] = 798;
        test_data[911] = 33'd8490724298;
        test_addr[912] = 238;
        test_data[912] = 33'd4586319590;
        test_addr[913] = 291;
        test_data[913] = 33'd3655503747;
        test_addr[914] = 329;
        test_data[914] = 33'd3903899561;
        test_addr[915] = 144;
        test_data[915] = 33'd4214779887;
        test_addr[916] = 691;
        test_data[916] = 33'd7121426868;
        test_addr[917] = 816;
        test_data[917] = 33'd912381185;
        test_addr[918] = 404;
        test_data[918] = 33'd4509066012;
        test_addr[919] = 541;
        test_data[919] = 33'd8503807599;
        test_addr[920] = 304;
        test_data[920] = 33'd3014575534;
        test_addr[921] = 108;
        test_data[921] = 33'd52659899;
        test_addr[922] = 932;
        test_data[922] = 33'd1290708529;
        test_addr[923] = 750;
        test_data[923] = 33'd380224476;
        test_addr[924] = 122;
        test_data[924] = 33'd1522076612;
        test_addr[925] = 845;
        test_data[925] = 33'd1963746399;
        test_addr[926] = 336;
        test_data[926] = 33'd6677673339;
        test_addr[927] = 658;
        test_data[927] = 33'd6371703314;
        test_addr[928] = 278;
        test_data[928] = 33'd3400886719;
        test_addr[929] = 531;
        test_data[929] = 33'd3479564107;
        test_addr[930] = 599;
        test_data[930] = 33'd7041741567;
        test_addr[931] = 978;
        test_data[931] = 33'd7873446819;
        test_addr[932] = 19;
        test_data[932] = 33'd2420327030;
        test_addr[933] = 196;
        test_data[933] = 33'd751103529;
        test_addr[934] = 427;
        test_data[934] = 33'd3998550133;
        test_addr[935] = 67;
        test_data[935] = 33'd3639768664;
        test_addr[936] = 319;
        test_data[936] = 33'd8248770922;
        test_addr[937] = 87;
        test_data[937] = 33'd8217428952;
        test_addr[938] = 1011;
        test_data[938] = 33'd2124493682;
        test_addr[939] = 74;
        test_data[939] = 33'd3405503829;
        test_addr[940] = 123;
        test_data[940] = 33'd3515538989;
        test_addr[941] = 421;
        test_data[941] = 33'd4143387137;
        test_addr[942] = 18;
        test_data[942] = 33'd3370794791;
        test_addr[943] = 10;
        test_data[943] = 33'd3594809116;
        test_addr[944] = 885;
        test_data[944] = 33'd728215166;
        test_addr[945] = 892;
        test_data[945] = 33'd7976219345;
        test_addr[946] = 879;
        test_data[946] = 33'd2227416794;
        test_addr[947] = 925;
        test_data[947] = 33'd1783235354;
        test_addr[948] = 967;
        test_data[948] = 33'd5738237391;
        test_addr[949] = 140;
        test_data[949] = 33'd3005608887;
        test_addr[950] = 166;
        test_data[950] = 33'd1217876369;
        test_addr[951] = 24;
        test_data[951] = 33'd1503049;
        test_addr[952] = 494;
        test_data[952] = 33'd1192454332;
        test_addr[953] = 457;
        test_data[953] = 33'd778796395;
        test_addr[954] = 61;
        test_data[954] = 33'd3243858099;
        test_addr[955] = 520;
        test_data[955] = 33'd3912596110;
        test_addr[956] = 414;
        test_data[956] = 33'd402300966;
        test_addr[957] = 0;
        test_data[957] = 33'd6235915199;
        test_addr[958] = 180;
        test_data[958] = 33'd4026446541;
        test_addr[959] = 708;
        test_data[959] = 33'd3363550927;
        test_addr[960] = 728;
        test_data[960] = 33'd6072302655;
        test_addr[961] = 655;
        test_data[961] = 33'd2678884701;
        test_addr[962] = 790;
        test_data[962] = 33'd5240800326;
        test_addr[963] = 116;
        test_data[963] = 33'd5752137139;
        test_addr[964] = 775;
        test_data[964] = 33'd4264175710;
        test_addr[965] = 39;
        test_data[965] = 33'd7929102593;
        test_addr[966] = 655;
        test_data[966] = 33'd2678884701;
        test_addr[967] = 924;
        test_data[967] = 33'd7156823247;
        test_addr[968] = 686;
        test_data[968] = 33'd318457616;
        test_addr[969] = 747;
        test_data[969] = 33'd4267106846;
        test_addr[970] = 585;
        test_data[970] = 33'd3586969900;
        test_addr[971] = 347;
        test_data[971] = 33'd8169775945;
        test_addr[972] = 909;
        test_data[972] = 33'd4367288555;
        test_addr[973] = 703;
        test_data[973] = 33'd7267050392;
        test_addr[974] = 923;
        test_data[974] = 33'd2479546912;
        test_addr[975] = 151;
        test_data[975] = 33'd5332051567;
        test_addr[976] = 681;
        test_data[976] = 33'd6006068068;
        test_addr[977] = 297;
        test_data[977] = 33'd7377276642;
        test_addr[978] = 255;
        test_data[978] = 33'd6211792075;
        test_addr[979] = 567;
        test_data[979] = 33'd806218001;
        test_addr[980] = 692;
        test_data[980] = 33'd4661411114;
        test_addr[981] = 869;
        test_data[981] = 33'd6631459962;
        test_addr[982] = 924;
        test_data[982] = 33'd7009780729;
        test_addr[983] = 833;
        test_data[983] = 33'd893301933;
        test_addr[984] = 1009;
        test_data[984] = 33'd2054454801;
        test_addr[985] = 997;
        test_data[985] = 33'd8276763053;
        test_addr[986] = 768;
        test_data[986] = 33'd3795726059;
        test_addr[987] = 346;
        test_data[987] = 33'd3114256567;
        test_addr[988] = 806;
        test_data[988] = 33'd7634373955;
        test_addr[989] = 378;
        test_data[989] = 33'd6762498788;
        test_addr[990] = 436;
        test_data[990] = 33'd1971182400;
        test_addr[991] = 467;
        test_data[991] = 33'd2928862965;
        test_addr[992] = 993;
        test_data[992] = 33'd2909818976;
        test_addr[993] = 852;
        test_data[993] = 33'd2596612030;
        test_addr[994] = 122;
        test_data[994] = 33'd1522076612;
        test_addr[995] = 964;
        test_data[995] = 33'd1077138145;
        test_addr[996] = 597;
        test_data[996] = 33'd572393240;
        test_addr[997] = 870;
        test_data[997] = 33'd166692004;
        test_addr[998] = 394;
        test_data[998] = 33'd5526543785;
        test_addr[999] = 344;
        test_data[999] = 33'd253890222;
        test_addr[1000] = 414;
        test_data[1000] = 33'd402300966;
        test_addr[1001] = 856;
        test_data[1001] = 33'd975862316;
        test_addr[1002] = 412;
        test_data[1002] = 33'd5982772419;
        test_addr[1003] = 71;
        test_data[1003] = 33'd3950328245;
        test_addr[1004] = 777;
        test_data[1004] = 33'd6001904970;
        test_addr[1005] = 907;
        test_data[1005] = 33'd4168846095;
        test_addr[1006] = 468;
        test_data[1006] = 33'd2002255513;
        test_addr[1007] = 721;
        test_data[1007] = 33'd8216915716;
        test_addr[1008] = 762;
        test_data[1008] = 33'd8542712035;
        test_addr[1009] = 107;
        test_data[1009] = 33'd4243198286;
        test_addr[1010] = 150;
        test_data[1010] = 33'd5030875849;
        test_addr[1011] = 719;
        test_data[1011] = 33'd3780764175;
        test_addr[1012] = 525;
        test_data[1012] = 33'd2628982812;
        test_addr[1013] = 566;
        test_data[1013] = 33'd770002620;
        test_addr[1014] = 286;
        test_data[1014] = 33'd2360048588;
        test_addr[1015] = 296;
        test_data[1015] = 33'd6676242800;
        test_addr[1016] = 868;
        test_data[1016] = 33'd2528507951;
        test_addr[1017] = 1015;
        test_data[1017] = 33'd2062647632;
        test_addr[1018] = 925;
        test_data[1018] = 33'd1783235354;
        test_addr[1019] = 931;
        test_data[1019] = 33'd2803979244;
        test_addr[1020] = 362;
        test_data[1020] = 33'd4225808861;
        test_addr[1021] = 917;
        test_data[1021] = 33'd6392673288;
        test_addr[1022] = 806;
        test_data[1022] = 33'd3339406659;
        test_addr[1023] = 628;
        test_data[1023] = 33'd7739780114;
        test_addr[1024] = 148;
        test_data[1024] = 33'd6194890702;
        test_addr[1025] = 651;
        test_data[1025] = 33'd1815633715;
        test_addr[1026] = 278;
        test_data[1026] = 33'd8148818173;
        test_addr[1027] = 632;
        test_data[1027] = 33'd162213990;
        test_addr[1028] = 552;
        test_data[1028] = 33'd6925457233;
        test_addr[1029] = 756;
        test_data[1029] = 33'd6387432324;
        test_addr[1030] = 296;
        test_data[1030] = 33'd2381275504;
        test_addr[1031] = 385;
        test_data[1031] = 33'd5417843210;
        test_addr[1032] = 184;
        test_data[1032] = 33'd3840564828;
        test_addr[1033] = 833;
        test_data[1033] = 33'd6186937878;
        test_addr[1034] = 746;
        test_data[1034] = 33'd2332255621;
        test_addr[1035] = 696;
        test_data[1035] = 33'd2694337344;
        test_addr[1036] = 202;
        test_data[1036] = 33'd5825244647;
        test_addr[1037] = 614;
        test_data[1037] = 33'd58076955;
        test_addr[1038] = 884;
        test_data[1038] = 33'd1323552558;
        test_addr[1039] = 977;
        test_data[1039] = 33'd1687923687;
        test_addr[1040] = 487;
        test_data[1040] = 33'd8185729776;
        test_addr[1041] = 401;
        test_data[1041] = 33'd7094310900;
        test_addr[1042] = 545;
        test_data[1042] = 33'd3465705991;
        test_addr[1043] = 7;
        test_data[1043] = 33'd7252660218;
        test_addr[1044] = 695;
        test_data[1044] = 33'd2186911345;
        test_addr[1045] = 559;
        test_data[1045] = 33'd7588610390;
        test_addr[1046] = 864;
        test_data[1046] = 33'd1571587926;
        test_addr[1047] = 972;
        test_data[1047] = 33'd3577819553;
        test_addr[1048] = 870;
        test_data[1048] = 33'd166692004;
        test_addr[1049] = 647;
        test_data[1049] = 33'd6946119;
        test_addr[1050] = 940;
        test_data[1050] = 33'd758677715;
        test_addr[1051] = 61;
        test_data[1051] = 33'd3243858099;
        test_addr[1052] = 140;
        test_data[1052] = 33'd7457150811;
        test_addr[1053] = 305;
        test_data[1053] = 33'd5396656275;
        test_addr[1054] = 258;
        test_data[1054] = 33'd2974304192;
        test_addr[1055] = 857;
        test_data[1055] = 33'd2261474441;
        test_addr[1056] = 307;
        test_data[1056] = 33'd6634543282;
        test_addr[1057] = 279;
        test_data[1057] = 33'd6144202271;
        test_addr[1058] = 855;
        test_data[1058] = 33'd6866220946;
        test_addr[1059] = 196;
        test_data[1059] = 33'd751103529;
        test_addr[1060] = 832;
        test_data[1060] = 33'd351971474;
        test_addr[1061] = 916;
        test_data[1061] = 33'd1736915697;
        test_addr[1062] = 948;
        test_data[1062] = 33'd716515165;
        test_addr[1063] = 865;
        test_data[1063] = 33'd1605398418;
        test_addr[1064] = 137;
        test_data[1064] = 33'd1215535519;
        test_addr[1065] = 970;
        test_data[1065] = 33'd1829669242;
        test_addr[1066] = 485;
        test_data[1066] = 33'd5495831061;
        test_addr[1067] = 747;
        test_data[1067] = 33'd4661830990;
        test_addr[1068] = 959;
        test_data[1068] = 33'd5205099699;
        test_addr[1069] = 290;
        test_data[1069] = 33'd3989670362;
        test_addr[1070] = 762;
        test_data[1070] = 33'd4247744739;
        test_addr[1071] = 83;
        test_data[1071] = 33'd5975311783;
        test_addr[1072] = 174;
        test_data[1072] = 33'd3604100316;
        test_addr[1073] = 590;
        test_data[1073] = 33'd1707606770;
        test_addr[1074] = 949;
        test_data[1074] = 33'd1458535013;
        test_addr[1075] = 638;
        test_data[1075] = 33'd2155582926;
        test_addr[1076] = 940;
        test_data[1076] = 33'd758677715;
        test_addr[1077] = 187;
        test_data[1077] = 33'd7297287928;
        test_addr[1078] = 54;
        test_data[1078] = 33'd2589183808;
        test_addr[1079] = 483;
        test_data[1079] = 33'd1178549137;
        test_addr[1080] = 478;
        test_data[1080] = 33'd627300334;
        test_addr[1081] = 159;
        test_data[1081] = 33'd4866761547;
        test_addr[1082] = 853;
        test_data[1082] = 33'd5783856874;
        test_addr[1083] = 831;
        test_data[1083] = 33'd992727670;
        test_addr[1084] = 727;
        test_data[1084] = 33'd2717525231;
        test_addr[1085] = 640;
        test_data[1085] = 33'd6017926257;
        test_addr[1086] = 4;
        test_data[1086] = 33'd1317783482;
        test_addr[1087] = 360;
        test_data[1087] = 33'd4335457434;
        test_addr[1088] = 312;
        test_data[1088] = 33'd1985873362;
        test_addr[1089] = 669;
        test_data[1089] = 33'd6798767308;
        test_addr[1090] = 717;
        test_data[1090] = 33'd2826264325;
        test_addr[1091] = 807;
        test_data[1091] = 33'd8440433509;
        test_addr[1092] = 733;
        test_data[1092] = 33'd7659479330;
        test_addr[1093] = 898;
        test_data[1093] = 33'd4064606830;
        test_addr[1094] = 846;
        test_data[1094] = 33'd2063463330;
        test_addr[1095] = 936;
        test_data[1095] = 33'd93762480;
        test_addr[1096] = 689;
        test_data[1096] = 33'd1681318426;
        test_addr[1097] = 775;
        test_data[1097] = 33'd4264175710;
        test_addr[1098] = 174;
        test_data[1098] = 33'd3604100316;
        test_addr[1099] = 415;
        test_data[1099] = 33'd5580768951;
        test_addr[1100] = 141;
        test_data[1100] = 33'd324907900;
        test_addr[1101] = 588;
        test_data[1101] = 33'd4041263385;
        test_addr[1102] = 848;
        test_data[1102] = 33'd1986134956;
        test_addr[1103] = 697;
        test_data[1103] = 33'd3089205481;
        test_addr[1104] = 160;
        test_data[1104] = 33'd5067522371;
        test_addr[1105] = 583;
        test_data[1105] = 33'd6183520255;
        test_addr[1106] = 1011;
        test_data[1106] = 33'd8290631108;
        test_addr[1107] = 749;
        test_data[1107] = 33'd1001567470;
        test_addr[1108] = 274;
        test_data[1108] = 33'd3318236443;
        test_addr[1109] = 340;
        test_data[1109] = 33'd3309872861;
        test_addr[1110] = 130;
        test_data[1110] = 33'd1268433295;
        test_addr[1111] = 557;
        test_data[1111] = 33'd4539639258;
        test_addr[1112] = 425;
        test_data[1112] = 33'd3540322948;
        test_addr[1113] = 204;
        test_data[1113] = 33'd5977734978;
        test_addr[1114] = 30;
        test_data[1114] = 33'd4880586894;
        test_addr[1115] = 982;
        test_data[1115] = 33'd772091063;
        test_addr[1116] = 975;
        test_data[1116] = 33'd1686953869;
        test_addr[1117] = 640;
        test_data[1117] = 33'd1722958961;
        test_addr[1118] = 761;
        test_data[1118] = 33'd2774007604;
        test_addr[1119] = 671;
        test_data[1119] = 33'd6965218581;
        test_addr[1120] = 853;
        test_data[1120] = 33'd7894501800;
        test_addr[1121] = 380;
        test_data[1121] = 33'd1024754085;
        test_addr[1122] = 717;
        test_data[1122] = 33'd6397259164;
        test_addr[1123] = 127;
        test_data[1123] = 33'd1731432911;
        test_addr[1124] = 668;
        test_data[1124] = 33'd977172141;
        test_addr[1125] = 376;
        test_data[1125] = 33'd3017136644;
        test_addr[1126] = 15;
        test_data[1126] = 33'd7484654752;
        test_addr[1127] = 619;
        test_data[1127] = 33'd1927924971;
        test_addr[1128] = 410;
        test_data[1128] = 33'd3405405453;
        test_addr[1129] = 873;
        test_data[1129] = 33'd722926779;
        test_addr[1130] = 841;
        test_data[1130] = 33'd124879403;
        test_addr[1131] = 911;
        test_data[1131] = 33'd6699783489;
        test_addr[1132] = 714;
        test_data[1132] = 33'd761390289;
        test_addr[1133] = 44;
        test_data[1133] = 33'd1301135708;
        test_addr[1134] = 512;
        test_data[1134] = 33'd112430786;
        test_addr[1135] = 672;
        test_data[1135] = 33'd3252626599;
        test_addr[1136] = 735;
        test_data[1136] = 33'd4187580926;
        test_addr[1137] = 318;
        test_data[1137] = 33'd1218864492;
        test_addr[1138] = 527;
        test_data[1138] = 33'd1169423377;
        test_addr[1139] = 1010;
        test_data[1139] = 33'd894431798;
        test_addr[1140] = 764;
        test_data[1140] = 33'd4377638901;
        test_addr[1141] = 524;
        test_data[1141] = 33'd6885604784;
        test_addr[1142] = 578;
        test_data[1142] = 33'd5557344247;
        test_addr[1143] = 647;
        test_data[1143] = 33'd5137056008;
        test_addr[1144] = 547;
        test_data[1144] = 33'd3100408585;
        test_addr[1145] = 429;
        test_data[1145] = 33'd6996815379;
        test_addr[1146] = 365;
        test_data[1146] = 33'd369210451;
        test_addr[1147] = 20;
        test_data[1147] = 33'd4648565853;
        test_addr[1148] = 509;
        test_data[1148] = 33'd1404134308;
        test_addr[1149] = 348;
        test_data[1149] = 33'd4786799480;
        test_addr[1150] = 490;
        test_data[1150] = 33'd755275238;
        test_addr[1151] = 196;
        test_data[1151] = 33'd751103529;
        test_addr[1152] = 113;
        test_data[1152] = 33'd2590394246;
        test_addr[1153] = 386;
        test_data[1153] = 33'd3669660999;
        test_addr[1154] = 339;
        test_data[1154] = 33'd4527677825;
        test_addr[1155] = 782;
        test_data[1155] = 33'd7722047099;
        test_addr[1156] = 843;
        test_data[1156] = 33'd7477027267;
        test_addr[1157] = 903;
        test_data[1157] = 33'd2634020074;
        test_addr[1158] = 35;
        test_data[1158] = 33'd1427007413;
        test_addr[1159] = 48;
        test_data[1159] = 33'd3748276960;
        test_addr[1160] = 981;
        test_data[1160] = 33'd5516712071;
        test_addr[1161] = 245;
        test_data[1161] = 33'd2052459312;
        test_addr[1162] = 589;
        test_data[1162] = 33'd1283209101;
        test_addr[1163] = 857;
        test_data[1163] = 33'd5613532770;
        test_addr[1164] = 486;
        test_data[1164] = 33'd2789818792;
        test_addr[1165] = 178;
        test_data[1165] = 33'd7204057384;
        test_addr[1166] = 254;
        test_data[1166] = 33'd4032840749;
        test_addr[1167] = 721;
        test_data[1167] = 33'd3921948420;
        test_addr[1168] = 606;
        test_data[1168] = 33'd4026351905;
        test_addr[1169] = 381;
        test_data[1169] = 33'd6133778541;
        test_addr[1170] = 182;
        test_data[1170] = 33'd2294431329;
        test_addr[1171] = 909;
        test_data[1171] = 33'd72321259;
        test_addr[1172] = 23;
        test_data[1172] = 33'd2154342992;
        test_addr[1173] = 827;
        test_data[1173] = 33'd4136395276;
        test_addr[1174] = 681;
        test_data[1174] = 33'd1711100772;
        test_addr[1175] = 111;
        test_data[1175] = 33'd3462749259;
        test_addr[1176] = 77;
        test_data[1176] = 33'd223605785;
        test_addr[1177] = 147;
        test_data[1177] = 33'd2764225137;
        test_addr[1178] = 344;
        test_data[1178] = 33'd253890222;
        test_addr[1179] = 674;
        test_data[1179] = 33'd2656360569;
        test_addr[1180] = 637;
        test_data[1180] = 33'd1672692856;
        test_addr[1181] = 761;
        test_data[1181] = 33'd2774007604;
        test_addr[1182] = 597;
        test_data[1182] = 33'd572393240;
        test_addr[1183] = 778;
        test_data[1183] = 33'd7509545295;
        test_addr[1184] = 807;
        test_data[1184] = 33'd4145466213;
        test_addr[1185] = 135;
        test_data[1185] = 33'd69857205;
        test_addr[1186] = 290;
        test_data[1186] = 33'd3989670362;
        test_addr[1187] = 735;
        test_data[1187] = 33'd4187580926;
        test_addr[1188] = 949;
        test_data[1188] = 33'd5933366934;
        test_addr[1189] = 487;
        test_data[1189] = 33'd5629918642;
        test_addr[1190] = 748;
        test_data[1190] = 33'd803782110;
        test_addr[1191] = 29;
        test_data[1191] = 33'd131073219;
        test_addr[1192] = 128;
        test_data[1192] = 33'd1320669106;
        test_addr[1193] = 791;
        test_data[1193] = 33'd6033689281;
        test_addr[1194] = 266;
        test_data[1194] = 33'd4857947400;
        test_addr[1195] = 96;
        test_data[1195] = 33'd7422710619;
        test_addr[1196] = 276;
        test_data[1196] = 33'd2694496543;
        test_addr[1197] = 417;
        test_data[1197] = 33'd2268883569;
        test_addr[1198] = 857;
        test_data[1198] = 33'd5747394507;
        test_addr[1199] = 356;
        test_data[1199] = 33'd4988367006;
        test_addr[1200] = 70;
        test_data[1200] = 33'd1368704711;
        test_addr[1201] = 186;
        test_data[1201] = 33'd275959827;
        test_addr[1202] = 191;
        test_data[1202] = 33'd4429539563;
        test_addr[1203] = 867;
        test_data[1203] = 33'd18555133;
        test_addr[1204] = 566;
        test_data[1204] = 33'd5659319685;
        test_addr[1205] = 386;
        test_data[1205] = 33'd3669660999;
        test_addr[1206] = 828;
        test_data[1206] = 33'd255493806;
        test_addr[1207] = 432;
        test_data[1207] = 33'd1268587008;
        test_addr[1208] = 948;
        test_data[1208] = 33'd716515165;
        test_addr[1209] = 621;
        test_data[1209] = 33'd1890719812;
        test_addr[1210] = 24;
        test_data[1210] = 33'd5645851620;
        test_addr[1211] = 165;
        test_data[1211] = 33'd106644142;
        test_addr[1212] = 780;
        test_data[1212] = 33'd404411201;
        test_addr[1213] = 620;
        test_data[1213] = 33'd3168866381;
        test_addr[1214] = 196;
        test_data[1214] = 33'd4513589842;
        test_addr[1215] = 647;
        test_data[1215] = 33'd842088712;
        test_addr[1216] = 966;
        test_data[1216] = 33'd1835137690;
        test_addr[1217] = 483;
        test_data[1217] = 33'd1178549137;
        test_addr[1218] = 113;
        test_data[1218] = 33'd2590394246;
        test_addr[1219] = 669;
        test_data[1219] = 33'd2503800012;
        test_addr[1220] = 435;
        test_data[1220] = 33'd3843532341;
        test_addr[1221] = 201;
        test_data[1221] = 33'd29735866;
        test_addr[1222] = 685;
        test_data[1222] = 33'd6708763506;
        test_addr[1223] = 667;
        test_data[1223] = 33'd3561967518;
        test_addr[1224] = 147;
        test_data[1224] = 33'd2764225137;
        test_addr[1225] = 97;
        test_data[1225] = 33'd5673895031;
        test_addr[1226] = 914;
        test_data[1226] = 33'd3697790821;
        test_addr[1227] = 206;
        test_data[1227] = 33'd380753888;
        test_addr[1228] = 63;
        test_data[1228] = 33'd6927994848;
        test_addr[1229] = 854;
        test_data[1229] = 33'd2260897852;
        test_addr[1230] = 474;
        test_data[1230] = 33'd4127845043;
        test_addr[1231] = 781;
        test_data[1231] = 33'd2061765198;
        test_addr[1232] = 349;
        test_data[1232] = 33'd7042377147;
        test_addr[1233] = 932;
        test_data[1233] = 33'd4657303822;
        test_addr[1234] = 491;
        test_data[1234] = 33'd2211071192;
        test_addr[1235] = 33;
        test_data[1235] = 33'd5779656203;
        test_addr[1236] = 218;
        test_data[1236] = 33'd4389591455;
        test_addr[1237] = 952;
        test_data[1237] = 33'd702855526;
        test_addr[1238] = 397;
        test_data[1238] = 33'd2491507040;
        test_addr[1239] = 700;
        test_data[1239] = 33'd759042820;
        test_addr[1240] = 564;
        test_data[1240] = 33'd7247987859;
        test_addr[1241] = 17;
        test_data[1241] = 33'd2023586953;
        test_addr[1242] = 640;
        test_data[1242] = 33'd6608778904;
        test_addr[1243] = 753;
        test_data[1243] = 33'd4949755487;
        test_addr[1244] = 501;
        test_data[1244] = 33'd7918829229;
        test_addr[1245] = 72;
        test_data[1245] = 33'd2563905635;
        test_addr[1246] = 596;
        test_data[1246] = 33'd4087896024;
        test_addr[1247] = 909;
        test_data[1247] = 33'd6544554853;
        test_addr[1248] = 717;
        test_data[1248] = 33'd2102291868;
        test_addr[1249] = 99;
        test_data[1249] = 33'd7175024271;
        test_addr[1250] = 11;
        test_data[1250] = 33'd3681162206;
        test_addr[1251] = 289;
        test_data[1251] = 33'd6326151339;
        test_addr[1252] = 262;
        test_data[1252] = 33'd4191130667;
        test_addr[1253] = 985;
        test_data[1253] = 33'd2974518957;
        test_addr[1254] = 89;
        test_data[1254] = 33'd3855383794;
        test_addr[1255] = 248;
        test_data[1255] = 33'd810408981;
        test_addr[1256] = 501;
        test_data[1256] = 33'd3623861933;
        test_addr[1257] = 64;
        test_data[1257] = 33'd3038722049;
        test_addr[1258] = 358;
        test_data[1258] = 33'd3979567529;
        test_addr[1259] = 355;
        test_data[1259] = 33'd3862589515;
        test_addr[1260] = 539;
        test_data[1260] = 33'd7702982231;
        test_addr[1261] = 310;
        test_data[1261] = 33'd3692301779;
        test_addr[1262] = 295;
        test_data[1262] = 33'd5377609965;
        test_addr[1263] = 784;
        test_data[1263] = 33'd4161914853;
        test_addr[1264] = 169;
        test_data[1264] = 33'd6111122785;
        test_addr[1265] = 927;
        test_data[1265] = 33'd1927721038;
        test_addr[1266] = 302;
        test_data[1266] = 33'd5057292467;
        test_addr[1267] = 179;
        test_data[1267] = 33'd3433493149;
        test_addr[1268] = 48;
        test_data[1268] = 33'd3748276960;
        test_addr[1269] = 756;
        test_data[1269] = 33'd2092465028;
        test_addr[1270] = 911;
        test_data[1270] = 33'd5832476673;
        test_addr[1271] = 209;
        test_data[1271] = 33'd6480062020;
        test_addr[1272] = 22;
        test_data[1272] = 33'd9397193;
        test_addr[1273] = 223;
        test_data[1273] = 33'd7818242704;
        test_addr[1274] = 712;
        test_data[1274] = 33'd1104352139;
        test_addr[1275] = 373;
        test_data[1275] = 33'd4405041255;
        test_addr[1276] = 314;
        test_data[1276] = 33'd751501571;
        test_addr[1277] = 909;
        test_data[1277] = 33'd2249587557;
        test_addr[1278] = 842;
        test_data[1278] = 33'd2581989200;
        test_addr[1279] = 922;
        test_data[1279] = 33'd715587172;
        test_addr[1280] = 954;
        test_data[1280] = 33'd5889637918;
        test_addr[1281] = 491;
        test_data[1281] = 33'd2211071192;
        test_addr[1282] = 677;
        test_data[1282] = 33'd4086784515;
        test_addr[1283] = 1000;
        test_data[1283] = 33'd5564630869;
        test_addr[1284] = 467;
        test_data[1284] = 33'd2928862965;
        test_addr[1285] = 77;
        test_data[1285] = 33'd223605785;
        test_addr[1286] = 773;
        test_data[1286] = 33'd1142927326;
        test_addr[1287] = 512;
        test_data[1287] = 33'd112430786;
        test_addr[1288] = 46;
        test_data[1288] = 33'd8390875893;
        test_addr[1289] = 344;
        test_data[1289] = 33'd253890222;
        test_addr[1290] = 348;
        test_data[1290] = 33'd7517394767;
        test_addr[1291] = 759;
        test_data[1291] = 33'd6483821833;
        test_addr[1292] = 840;
        test_data[1292] = 33'd5083816483;
        test_addr[1293] = 315;
        test_data[1293] = 33'd7872459330;
        test_addr[1294] = 766;
        test_data[1294] = 33'd6099268808;
        test_addr[1295] = 660;
        test_data[1295] = 33'd6121690392;
        test_addr[1296] = 542;
        test_data[1296] = 33'd6983338126;
        test_addr[1297] = 696;
        test_data[1297] = 33'd2694337344;
        test_addr[1298] = 731;
        test_data[1298] = 33'd1134545885;
        test_addr[1299] = 588;
        test_data[1299] = 33'd4041263385;
        test_addr[1300] = 218;
        test_data[1300] = 33'd94624159;
        test_addr[1301] = 815;
        test_data[1301] = 33'd1640602374;
        test_addr[1302] = 981;
        test_data[1302] = 33'd1221744775;
        test_addr[1303] = 852;
        test_data[1303] = 33'd7272401185;
        test_addr[1304] = 895;
        test_data[1304] = 33'd2540543346;
        test_addr[1305] = 538;
        test_data[1305] = 33'd1157057488;
        test_addr[1306] = 242;
        test_data[1306] = 33'd1982815146;
        test_addr[1307] = 717;
        test_data[1307] = 33'd2102291868;
        test_addr[1308] = 594;
        test_data[1308] = 33'd3790697293;
        test_addr[1309] = 462;
        test_data[1309] = 33'd8164776817;
        test_addr[1310] = 223;
        test_data[1310] = 33'd7505045586;
        test_addr[1311] = 463;
        test_data[1311] = 33'd1603013143;
        test_addr[1312] = 1007;
        test_data[1312] = 33'd3354638094;
        test_addr[1313] = 376;
        test_data[1313] = 33'd3017136644;
        test_addr[1314] = 41;
        test_data[1314] = 33'd6033521857;
        test_addr[1315] = 604;
        test_data[1315] = 33'd70723367;
        test_addr[1316] = 54;
        test_data[1316] = 33'd8562339813;
        test_addr[1317] = 184;
        test_data[1317] = 33'd3840564828;
        test_addr[1318] = 847;
        test_data[1318] = 33'd196428976;
        test_addr[1319] = 69;
        test_data[1319] = 33'd1753936223;
        test_addr[1320] = 232;
        test_data[1320] = 33'd930589679;
        test_addr[1321] = 828;
        test_data[1321] = 33'd6641429838;
        test_addr[1322] = 45;
        test_data[1322] = 33'd8056951560;
        test_addr[1323] = 219;
        test_data[1323] = 33'd308900539;
        test_addr[1324] = 663;
        test_data[1324] = 33'd1455377357;
        test_addr[1325] = 669;
        test_data[1325] = 33'd2503800012;
        test_addr[1326] = 119;
        test_data[1326] = 33'd2763234325;
        test_addr[1327] = 688;
        test_data[1327] = 33'd4133517367;
        test_addr[1328] = 297;
        test_data[1328] = 33'd3082309346;
        test_addr[1329] = 565;
        test_data[1329] = 33'd2843637762;
        test_addr[1330] = 780;
        test_data[1330] = 33'd404411201;
        test_addr[1331] = 571;
        test_data[1331] = 33'd3849053210;
        test_addr[1332] = 758;
        test_data[1332] = 33'd7660653570;
        test_addr[1333] = 470;
        test_data[1333] = 33'd4703955904;
        test_addr[1334] = 520;
        test_data[1334] = 33'd6944688602;
        test_addr[1335] = 931;
        test_data[1335] = 33'd2803979244;
        test_addr[1336] = 902;
        test_data[1336] = 33'd5709445376;
        test_addr[1337] = 911;
        test_data[1337] = 33'd1537509377;
        test_addr[1338] = 799;
        test_data[1338] = 33'd3954575845;
        test_addr[1339] = 870;
        test_data[1339] = 33'd166692004;
        test_addr[1340] = 106;
        test_data[1340] = 33'd898134430;
        test_addr[1341] = 339;
        test_data[1341] = 33'd232710529;
        test_addr[1342] = 356;
        test_data[1342] = 33'd6672956910;
        test_addr[1343] = 683;
        test_data[1343] = 33'd5392604401;
        test_addr[1344] = 658;
        test_data[1344] = 33'd2076736018;
        test_addr[1345] = 703;
        test_data[1345] = 33'd5209880850;
        test_addr[1346] = 979;
        test_data[1346] = 33'd1509757740;
        test_addr[1347] = 693;
        test_data[1347] = 33'd2069998988;
        test_addr[1348] = 23;
        test_data[1348] = 33'd2154342992;
        test_addr[1349] = 495;
        test_data[1349] = 33'd885613252;
        test_addr[1350] = 934;
        test_data[1350] = 33'd2539789535;
        test_addr[1351] = 912;
        test_data[1351] = 33'd1978461553;
        test_addr[1352] = 1007;
        test_data[1352] = 33'd3354638094;
        test_addr[1353] = 704;
        test_data[1353] = 33'd2320769301;
        test_addr[1354] = 357;
        test_data[1354] = 33'd4022908127;
        test_addr[1355] = 370;
        test_data[1355] = 33'd4551654172;
        test_addr[1356] = 154;
        test_data[1356] = 33'd6560321906;
        test_addr[1357] = 252;
        test_data[1357] = 33'd5468455138;
        test_addr[1358] = 303;
        test_data[1358] = 33'd6347969693;
        test_addr[1359] = 419;
        test_data[1359] = 33'd4133168253;
        test_addr[1360] = 102;
        test_data[1360] = 33'd1124317209;
        test_addr[1361] = 894;
        test_data[1361] = 33'd5516969405;
        test_addr[1362] = 37;
        test_data[1362] = 33'd4017425673;
        test_addr[1363] = 54;
        test_data[1363] = 33'd4853967616;
        test_addr[1364] = 1003;
        test_data[1364] = 33'd8442982682;
        test_addr[1365] = 131;
        test_data[1365] = 33'd813280569;
        test_addr[1366] = 730;
        test_data[1366] = 33'd2774040910;
        test_addr[1367] = 566;
        test_data[1367] = 33'd1364352389;
        test_addr[1368] = 260;
        test_data[1368] = 33'd3363163059;
        test_addr[1369] = 907;
        test_data[1369] = 33'd4168846095;
        test_addr[1370] = 578;
        test_data[1370] = 33'd1262376951;
        test_addr[1371] = 299;
        test_data[1371] = 33'd3707209855;
        test_addr[1372] = 602;
        test_data[1372] = 33'd7776071822;
        test_addr[1373] = 880;
        test_data[1373] = 33'd6419643479;
        test_addr[1374] = 109;
        test_data[1374] = 33'd2394762171;
        test_addr[1375] = 850;
        test_data[1375] = 33'd640217809;
        test_addr[1376] = 133;
        test_data[1376] = 33'd1645346336;
        test_addr[1377] = 927;
        test_data[1377] = 33'd1927721038;
        test_addr[1378] = 516;
        test_data[1378] = 33'd7530390101;
        test_addr[1379] = 257;
        test_data[1379] = 33'd7053270609;
        test_addr[1380] = 476;
        test_data[1380] = 33'd3010424531;
        test_addr[1381] = 330;
        test_data[1381] = 33'd7594307275;
        test_addr[1382] = 501;
        test_data[1382] = 33'd3623861933;
        test_addr[1383] = 638;
        test_data[1383] = 33'd2155582926;
        test_addr[1384] = 1017;
        test_data[1384] = 33'd5190891398;
        test_addr[1385] = 27;
        test_data[1385] = 33'd6617680999;
        test_addr[1386] = 802;
        test_data[1386] = 33'd8473857808;
        test_addr[1387] = 690;
        test_data[1387] = 33'd4095690594;
        test_addr[1388] = 1005;
        test_data[1388] = 33'd1098300837;
        test_addr[1389] = 343;
        test_data[1389] = 33'd2472167151;
        test_addr[1390] = 564;
        test_data[1390] = 33'd2953020563;
        test_addr[1391] = 317;
        test_data[1391] = 33'd7974375809;
        test_addr[1392] = 187;
        test_data[1392] = 33'd3002320632;
        test_addr[1393] = 280;
        test_data[1393] = 33'd5744733524;
        test_addr[1394] = 900;
        test_data[1394] = 33'd3715729542;
        test_addr[1395] = 251;
        test_data[1395] = 33'd5563861074;
        test_addr[1396] = 894;
        test_data[1396] = 33'd1222002109;
        test_addr[1397] = 515;
        test_data[1397] = 33'd1989592525;
        test_addr[1398] = 603;
        test_data[1398] = 33'd2447831809;
        test_addr[1399] = 186;
        test_data[1399] = 33'd5965245879;
        test_addr[1400] = 140;
        test_data[1400] = 33'd3162183515;
        test_addr[1401] = 834;
        test_data[1401] = 33'd5447660091;
        test_addr[1402] = 330;
        test_data[1402] = 33'd6357429645;
        test_addr[1403] = 278;
        test_data[1403] = 33'd3853850877;
        test_addr[1404] = 166;
        test_data[1404] = 33'd1217876369;
        test_addr[1405] = 61;
        test_data[1405] = 33'd3243858099;
        test_addr[1406] = 60;
        test_data[1406] = 33'd2895705112;
        test_addr[1407] = 1;
        test_data[1407] = 33'd2545176946;
        test_addr[1408] = 418;
        test_data[1408] = 33'd564521412;
        test_addr[1409] = 955;
        test_data[1409] = 33'd4217331207;
        test_addr[1410] = 199;
        test_data[1410] = 33'd6262982402;
        test_addr[1411] = 534;
        test_data[1411] = 33'd2464887914;
        test_addr[1412] = 940;
        test_data[1412] = 33'd7152119175;
        test_addr[1413] = 503;
        test_data[1413] = 33'd2825090233;
        test_addr[1414] = 940;
        test_data[1414] = 33'd2857151879;
        test_addr[1415] = 222;
        test_data[1415] = 33'd1146860549;
        test_addr[1416] = 554;
        test_data[1416] = 33'd2207183766;
        test_addr[1417] = 115;
        test_data[1417] = 33'd2347364473;
        test_addr[1418] = 714;
        test_data[1418] = 33'd761390289;
        test_addr[1419] = 273;
        test_data[1419] = 33'd56693191;
        test_addr[1420] = 70;
        test_data[1420] = 33'd1368704711;
        test_addr[1421] = 770;
        test_data[1421] = 33'd7548571949;
        test_addr[1422] = 939;
        test_data[1422] = 33'd536731119;
        test_addr[1423] = 321;
        test_data[1423] = 33'd6925867570;
        test_addr[1424] = 806;
        test_data[1424] = 33'd3339406659;
        test_addr[1425] = 833;
        test_data[1425] = 33'd1891970582;
        test_addr[1426] = 408;
        test_data[1426] = 33'd1130836166;
        test_addr[1427] = 472;
        test_data[1427] = 33'd2925733218;
        test_addr[1428] = 198;
        test_data[1428] = 33'd5896591301;
        test_addr[1429] = 321;
        test_data[1429] = 33'd2630900274;
        test_addr[1430] = 893;
        test_data[1430] = 33'd6228356496;
        test_addr[1431] = 365;
        test_data[1431] = 33'd369210451;
        test_addr[1432] = 590;
        test_data[1432] = 33'd1707606770;
        test_addr[1433] = 735;
        test_data[1433] = 33'd5523494548;
        test_addr[1434] = 851;
        test_data[1434] = 33'd550630034;
        test_addr[1435] = 87;
        test_data[1435] = 33'd3922461656;
        test_addr[1436] = 898;
        test_data[1436] = 33'd4064606830;
        test_addr[1437] = 405;
        test_data[1437] = 33'd516109638;
        test_addr[1438] = 377;
        test_data[1438] = 33'd2370864657;
        test_addr[1439] = 806;
        test_data[1439] = 33'd3339406659;
        test_addr[1440] = 973;
        test_data[1440] = 33'd5281772514;
        test_addr[1441] = 733;
        test_data[1441] = 33'd8005248793;
        test_addr[1442] = 617;
        test_data[1442] = 33'd6915372624;
        test_addr[1443] = 274;
        test_data[1443] = 33'd4485408491;
        test_addr[1444] = 908;
        test_data[1444] = 33'd1134632579;
        test_addr[1445] = 760;
        test_data[1445] = 33'd4199067864;
        test_addr[1446] = 446;
        test_data[1446] = 33'd6204434912;
        test_addr[1447] = 984;
        test_data[1447] = 33'd7463567831;
        test_addr[1448] = 40;
        test_data[1448] = 33'd2224301287;
        test_addr[1449] = 456;
        test_data[1449] = 33'd3608555727;
        test_addr[1450] = 492;
        test_data[1450] = 33'd2984910114;
        test_addr[1451] = 614;
        test_data[1451] = 33'd58076955;
        test_addr[1452] = 330;
        test_data[1452] = 33'd5720018780;
        test_addr[1453] = 329;
        test_data[1453] = 33'd3903899561;
        test_addr[1454] = 205;
        test_data[1454] = 33'd2173752367;
        test_addr[1455] = 260;
        test_data[1455] = 33'd3363163059;
        test_addr[1456] = 912;
        test_data[1456] = 33'd1978461553;
        test_addr[1457] = 621;
        test_data[1457] = 33'd1890719812;
        test_addr[1458] = 743;
        test_data[1458] = 33'd7907303613;
        test_addr[1459] = 895;
        test_data[1459] = 33'd6632829968;
        test_addr[1460] = 965;
        test_data[1460] = 33'd4354858199;
        test_addr[1461] = 768;
        test_data[1461] = 33'd3795726059;
        test_addr[1462] = 170;
        test_data[1462] = 33'd2103127943;
        test_addr[1463] = 976;
        test_data[1463] = 33'd3839524366;
        test_addr[1464] = 493;
        test_data[1464] = 33'd392841551;
        test_addr[1465] = 488;
        test_data[1465] = 33'd2484186896;
        test_addr[1466] = 532;
        test_data[1466] = 33'd7481466375;
        test_addr[1467] = 648;
        test_data[1467] = 33'd2025862340;
        test_addr[1468] = 695;
        test_data[1468] = 33'd2186911345;
        test_addr[1469] = 277;
        test_data[1469] = 33'd2799792130;
        test_addr[1470] = 624;
        test_data[1470] = 33'd8071541066;
        test_addr[1471] = 427;
        test_data[1471] = 33'd3998550133;
        test_addr[1472] = 719;
        test_data[1472] = 33'd3780764175;
        test_addr[1473] = 367;
        test_data[1473] = 33'd7047582222;
        test_addr[1474] = 113;
        test_data[1474] = 33'd6324911211;
        test_addr[1475] = 197;
        test_data[1475] = 33'd2393364357;
        test_addr[1476] = 590;
        test_data[1476] = 33'd4549509652;
        test_addr[1477] = 978;
        test_data[1477] = 33'd5904384292;
        test_addr[1478] = 948;
        test_data[1478] = 33'd6051245577;
        test_addr[1479] = 614;
        test_data[1479] = 33'd58076955;
        test_addr[1480] = 692;
        test_data[1480] = 33'd366443818;
        test_addr[1481] = 47;
        test_data[1481] = 33'd5979200969;
        test_addr[1482] = 221;
        test_data[1482] = 33'd720358563;
        test_addr[1483] = 762;
        test_data[1483] = 33'd4247744739;
        test_addr[1484] = 504;
        test_data[1484] = 33'd2373341895;
        test_addr[1485] = 858;
        test_data[1485] = 33'd5320593016;
        test_addr[1486] = 206;
        test_data[1486] = 33'd380753888;
        test_addr[1487] = 151;
        test_data[1487] = 33'd1037084271;
        test_addr[1488] = 453;
        test_data[1488] = 33'd3723143858;
        test_addr[1489] = 278;
        test_data[1489] = 33'd3853850877;
        test_addr[1490] = 274;
        test_data[1490] = 33'd190441195;
        test_addr[1491] = 668;
        test_data[1491] = 33'd977172141;
        test_addr[1492] = 984;
        test_data[1492] = 33'd3168600535;
        test_addr[1493] = 151;
        test_data[1493] = 33'd6421446107;
        test_addr[1494] = 938;
        test_data[1494] = 33'd1559360487;
        test_addr[1495] = 837;
        test_data[1495] = 33'd7042841169;
        test_addr[1496] = 192;
        test_data[1496] = 33'd2694434016;
        test_addr[1497] = 911;
        test_data[1497] = 33'd6342066238;
        test_addr[1498] = 699;
        test_data[1498] = 33'd6263778256;
        test_addr[1499] = 537;
        test_data[1499] = 33'd810473933;
        test_addr[1500] = 200;
        test_data[1500] = 33'd4007449550;
        test_addr[1501] = 425;
        test_data[1501] = 33'd3540322948;
        test_addr[1502] = 201;
        test_data[1502] = 33'd29735866;
        test_addr[1503] = 863;
        test_data[1503] = 33'd1325550564;
        test_addr[1504] = 204;
        test_data[1504] = 33'd1682767682;
        test_addr[1505] = 588;
        test_data[1505] = 33'd4041263385;
        test_addr[1506] = 696;
        test_data[1506] = 33'd2694337344;
        test_addr[1507] = 112;
        test_data[1507] = 33'd5585309931;
        test_addr[1508] = 179;
        test_data[1508] = 33'd3433493149;
        test_addr[1509] = 687;
        test_data[1509] = 33'd1000461927;
        test_addr[1510] = 766;
        test_data[1510] = 33'd1804301512;
        test_addr[1511] = 189;
        test_data[1511] = 33'd3994613051;
        test_addr[1512] = 21;
        test_data[1512] = 33'd1714185095;
        test_addr[1513] = 84;
        test_data[1513] = 33'd5189128390;
        test_addr[1514] = 129;
        test_data[1514] = 33'd1882082764;
        test_addr[1515] = 169;
        test_data[1515] = 33'd1816155489;
        test_addr[1516] = 138;
        test_data[1516] = 33'd2910298998;
        test_addr[1517] = 907;
        test_data[1517] = 33'd4168846095;
        test_addr[1518] = 115;
        test_data[1518] = 33'd2347364473;
        test_addr[1519] = 782;
        test_data[1519] = 33'd5067651649;
        test_addr[1520] = 252;
        test_data[1520] = 33'd1173487842;
        test_addr[1521] = 670;
        test_data[1521] = 33'd5908370301;
        test_addr[1522] = 909;
        test_data[1522] = 33'd8230962327;
        test_addr[1523] = 474;
        test_data[1523] = 33'd4127845043;
        test_addr[1524] = 477;
        test_data[1524] = 33'd2823642870;
        test_addr[1525] = 86;
        test_data[1525] = 33'd2898065894;
        test_addr[1526] = 221;
        test_data[1526] = 33'd720358563;
        test_addr[1527] = 506;
        test_data[1527] = 33'd7440261146;
        test_addr[1528] = 150;
        test_data[1528] = 33'd735908553;
        test_addr[1529] = 578;
        test_data[1529] = 33'd1262376951;
        test_addr[1530] = 392;
        test_data[1530] = 33'd6926277069;
        test_addr[1531] = 989;
        test_data[1531] = 33'd7107439867;
        test_addr[1532] = 776;
        test_data[1532] = 33'd769284591;
        test_addr[1533] = 218;
        test_data[1533] = 33'd94624159;
        test_addr[1534] = 556;
        test_data[1534] = 33'd2030797940;
        test_addr[1535] = 173;
        test_data[1535] = 33'd1456155483;
        test_addr[1536] = 905;
        test_data[1536] = 33'd3362997925;
        test_addr[1537] = 836;
        test_data[1537] = 33'd1052769268;
        test_addr[1538] = 509;
        test_data[1538] = 33'd8084294061;
        test_addr[1539] = 65;
        test_data[1539] = 33'd7233181161;
        test_addr[1540] = 53;
        test_data[1540] = 33'd421375381;
        test_addr[1541] = 142;
        test_data[1541] = 33'd2983160463;
        test_addr[1542] = 962;
        test_data[1542] = 33'd3905065194;
        test_addr[1543] = 245;
        test_data[1543] = 33'd2052459312;
        test_addr[1544] = 69;
        test_data[1544] = 33'd7202947070;
        test_addr[1545] = 826;
        test_data[1545] = 33'd690145171;
        test_addr[1546] = 580;
        test_data[1546] = 33'd436662051;
        test_addr[1547] = 317;
        test_data[1547] = 33'd7030568912;
        test_addr[1548] = 136;
        test_data[1548] = 33'd7314443525;
        test_addr[1549] = 846;
        test_data[1549] = 33'd5471318843;
        test_addr[1550] = 960;
        test_data[1550] = 33'd1495890564;
        test_addr[1551] = 106;
        test_data[1551] = 33'd898134430;
        test_addr[1552] = 20;
        test_data[1552] = 33'd8517755671;
        test_addr[1553] = 1007;
        test_data[1553] = 33'd3354638094;
        test_addr[1554] = 894;
        test_data[1554] = 33'd7074639747;
        test_addr[1555] = 584;
        test_data[1555] = 33'd3681182924;
        test_addr[1556] = 524;
        test_data[1556] = 33'd2590637488;
        test_addr[1557] = 822;
        test_data[1557] = 33'd534736813;
        test_addr[1558] = 634;
        test_data[1558] = 33'd2731773946;
        test_addr[1559] = 384;
        test_data[1559] = 33'd6072368523;
        test_addr[1560] = 727;
        test_data[1560] = 33'd2717525231;
        test_addr[1561] = 304;
        test_data[1561] = 33'd3014575534;
        test_addr[1562] = 592;
        test_data[1562] = 33'd938793682;
        test_addr[1563] = 651;
        test_data[1563] = 33'd5654066229;
        test_addr[1564] = 266;
        test_data[1564] = 33'd562980104;
        test_addr[1565] = 794;
        test_data[1565] = 33'd1458211943;
        test_addr[1566] = 159;
        test_data[1566] = 33'd571794251;
        test_addr[1567] = 324;
        test_data[1567] = 33'd330852185;
        test_addr[1568] = 91;
        test_data[1568] = 33'd3196504029;
        test_addr[1569] = 576;
        test_data[1569] = 33'd4983033453;
        test_addr[1570] = 446;
        test_data[1570] = 33'd1909467616;
        test_addr[1571] = 229;
        test_data[1571] = 33'd920626449;
        test_addr[1572] = 396;
        test_data[1572] = 33'd5234684424;
        test_addr[1573] = 542;
        test_data[1573] = 33'd2688370830;
        test_addr[1574] = 396;
        test_data[1574] = 33'd939717128;
        test_addr[1575] = 262;
        test_data[1575] = 33'd8260972120;
        test_addr[1576] = 253;
        test_data[1576] = 33'd2796634323;
        test_addr[1577] = 728;
        test_data[1577] = 33'd5101551394;
        test_addr[1578] = 436;
        test_data[1578] = 33'd1971182400;
        test_addr[1579] = 661;
        test_data[1579] = 33'd981018742;
        test_addr[1580] = 446;
        test_data[1580] = 33'd1909467616;
        test_addr[1581] = 27;
        test_data[1581] = 33'd2322713703;
        test_addr[1582] = 905;
        test_data[1582] = 33'd6967385077;
        test_addr[1583] = 23;
        test_data[1583] = 33'd5382366738;
        test_addr[1584] = 226;
        test_data[1584] = 33'd4004290607;
        test_addr[1585] = 550;
        test_data[1585] = 33'd2861464618;
        test_addr[1586] = 97;
        test_data[1586] = 33'd1378927735;
        test_addr[1587] = 36;
        test_data[1587] = 33'd7309348142;
        test_addr[1588] = 7;
        test_data[1588] = 33'd2957692922;
        test_addr[1589] = 324;
        test_data[1589] = 33'd330852185;
        test_addr[1590] = 997;
        test_data[1590] = 33'd3981795757;
        test_addr[1591] = 243;
        test_data[1591] = 33'd3048963064;
        test_addr[1592] = 442;
        test_data[1592] = 33'd1682936301;
        test_addr[1593] = 468;
        test_data[1593] = 33'd4344805153;
        test_addr[1594] = 819;
        test_data[1594] = 33'd7115811212;
        test_addr[1595] = 967;
        test_data[1595] = 33'd1443270095;
        test_addr[1596] = 972;
        test_data[1596] = 33'd7428902819;
        test_addr[1597] = 161;
        test_data[1597] = 33'd3641808353;
        test_addr[1598] = 93;
        test_data[1598] = 33'd263550839;
        test_addr[1599] = 9;
        test_data[1599] = 33'd7260278852;
        test_addr[1600] = 938;
        test_data[1600] = 33'd1559360487;
        test_addr[1601] = 621;
        test_data[1601] = 33'd1890719812;
        test_addr[1602] = 980;
        test_data[1602] = 33'd7889910182;
        test_addr[1603] = 1017;
        test_data[1603] = 33'd8010623804;
        test_addr[1604] = 997;
        test_data[1604] = 33'd3981795757;
        test_addr[1605] = 662;
        test_data[1605] = 33'd2183779360;
        test_addr[1606] = 910;
        test_data[1606] = 33'd5288809774;
        test_addr[1607] = 751;
        test_data[1607] = 33'd2723074538;
        test_addr[1608] = 204;
        test_data[1608] = 33'd1682767682;
        test_addr[1609] = 540;
        test_data[1609] = 33'd432267239;
        test_addr[1610] = 603;
        test_data[1610] = 33'd2447831809;
        test_addr[1611] = 1021;
        test_data[1611] = 33'd5688874170;
        test_addr[1612] = 437;
        test_data[1612] = 33'd3188866646;
        test_addr[1613] = 99;
        test_data[1613] = 33'd2880056975;
        test_addr[1614] = 429;
        test_data[1614] = 33'd2701848083;
        test_addr[1615] = 90;
        test_data[1615] = 33'd4119473539;
        test_addr[1616] = 389;
        test_data[1616] = 33'd2549642068;
        test_addr[1617] = 630;
        test_data[1617] = 33'd4437589608;
        test_addr[1618] = 345;
        test_data[1618] = 33'd2662284645;
        test_addr[1619] = 886;
        test_data[1619] = 33'd4267669502;
        test_addr[1620] = 740;
        test_data[1620] = 33'd6085180590;
        test_addr[1621] = 347;
        test_data[1621] = 33'd3874808649;
        test_addr[1622] = 331;
        test_data[1622] = 33'd3237563871;
        test_addr[1623] = 1018;
        test_data[1623] = 33'd7026150185;
        test_addr[1624] = 627;
        test_data[1624] = 33'd1310702174;
        test_addr[1625] = 849;
        test_data[1625] = 33'd1321707081;
        test_addr[1626] = 494;
        test_data[1626] = 33'd1192454332;
        test_addr[1627] = 157;
        test_data[1627] = 33'd6113838378;
        test_addr[1628] = 506;
        test_data[1628] = 33'd3145293850;
        test_addr[1629] = 702;
        test_data[1629] = 33'd7540665453;
        test_addr[1630] = 744;
        test_data[1630] = 33'd7099226051;
        test_addr[1631] = 59;
        test_data[1631] = 33'd7726204500;
        test_addr[1632] = 688;
        test_data[1632] = 33'd7297035982;
        test_addr[1633] = 298;
        test_data[1633] = 33'd1530159267;
        test_addr[1634] = 34;
        test_data[1634] = 33'd2988630753;
        test_addr[1635] = 335;
        test_data[1635] = 33'd6376729352;
        test_addr[1636] = 871;
        test_data[1636] = 33'd3900374916;
        test_addr[1637] = 716;
        test_data[1637] = 33'd1341092090;
        test_addr[1638] = 644;
        test_data[1638] = 33'd8105631119;
        test_addr[1639] = 772;
        test_data[1639] = 33'd3678900751;
        test_addr[1640] = 583;
        test_data[1640] = 33'd1888552959;
        test_addr[1641] = 559;
        test_data[1641] = 33'd3293643094;
        test_addr[1642] = 54;
        test_data[1642] = 33'd559000320;
        test_addr[1643] = 43;
        test_data[1643] = 33'd2636643983;
        test_addr[1644] = 653;
        test_data[1644] = 33'd6114678215;
        test_addr[1645] = 290;
        test_data[1645] = 33'd3989670362;
        test_addr[1646] = 37;
        test_data[1646] = 33'd7150942120;
        test_addr[1647] = 625;
        test_data[1647] = 33'd4643152190;
        test_addr[1648] = 179;
        test_data[1648] = 33'd3433493149;
        test_addr[1649] = 716;
        test_data[1649] = 33'd1341092090;
        test_addr[1650] = 131;
        test_data[1650] = 33'd813280569;
        test_addr[1651] = 523;
        test_data[1651] = 33'd577685601;
        test_addr[1652] = 504;
        test_data[1652] = 33'd2373341895;
        test_addr[1653] = 820;
        test_data[1653] = 33'd4175331955;
        test_addr[1654] = 214;
        test_data[1654] = 33'd3250589043;
        test_addr[1655] = 0;
        test_data[1655] = 33'd1940947903;
        test_addr[1656] = 835;
        test_data[1656] = 33'd3461985819;
        test_addr[1657] = 773;
        test_data[1657] = 33'd1142927326;
        test_addr[1658] = 145;
        test_data[1658] = 33'd1207656834;
        test_addr[1659] = 130;
        test_data[1659] = 33'd1268433295;
        test_addr[1660] = 703;
        test_data[1660] = 33'd4671088680;
        test_addr[1661] = 165;
        test_data[1661] = 33'd106644142;
        test_addr[1662] = 352;
        test_data[1662] = 33'd3944142242;
        test_addr[1663] = 916;
        test_data[1663] = 33'd1736915697;
        test_addr[1664] = 371;
        test_data[1664] = 33'd941454407;
        test_addr[1665] = 549;
        test_data[1665] = 33'd3755325729;
        test_addr[1666] = 848;
        test_data[1666] = 33'd1986134956;
        test_addr[1667] = 92;
        test_data[1667] = 33'd5525490977;
        test_addr[1668] = 94;
        test_data[1668] = 33'd2491615377;
        test_addr[1669] = 955;
        test_data[1669] = 33'd4494798025;
        test_addr[1670] = 270;
        test_data[1670] = 33'd2409706630;
        test_addr[1671] = 363;
        test_data[1671] = 33'd5688413322;
        test_addr[1672] = 466;
        test_data[1672] = 33'd633115602;
        test_addr[1673] = 227;
        test_data[1673] = 33'd905576619;
        test_addr[1674] = 661;
        test_data[1674] = 33'd981018742;
        test_addr[1675] = 103;
        test_data[1675] = 33'd4690276874;
        test_addr[1676] = 119;
        test_data[1676] = 33'd2763234325;
        test_addr[1677] = 783;
        test_data[1677] = 33'd2573492496;
        test_addr[1678] = 1015;
        test_data[1678] = 33'd2062647632;
        test_addr[1679] = 70;
        test_data[1679] = 33'd1368704711;
        test_addr[1680] = 489;
        test_data[1680] = 33'd7898133209;
        test_addr[1681] = 259;
        test_data[1681] = 33'd3390847646;
        test_addr[1682] = 282;
        test_data[1682] = 33'd5567263460;
        test_addr[1683] = 395;
        test_data[1683] = 33'd1292390397;
        test_addr[1684] = 874;
        test_data[1684] = 33'd2931664417;
        test_addr[1685] = 599;
        test_data[1685] = 33'd7154998828;
        test_addr[1686] = 188;
        test_data[1686] = 33'd4083814239;
        test_addr[1687] = 104;
        test_data[1687] = 33'd3714367826;
        test_addr[1688] = 598;
        test_data[1688] = 33'd3684002157;
        test_addr[1689] = 672;
        test_data[1689] = 33'd7590013900;
        test_addr[1690] = 269;
        test_data[1690] = 33'd2017951304;
        test_addr[1691] = 402;
        test_data[1691] = 33'd1208032225;
        test_addr[1692] = 707;
        test_data[1692] = 33'd5161085458;
        test_addr[1693] = 761;
        test_data[1693] = 33'd5255246887;
        test_addr[1694] = 570;
        test_data[1694] = 33'd1501919528;
        test_addr[1695] = 706;
        test_data[1695] = 33'd785242298;
        test_addr[1696] = 559;
        test_data[1696] = 33'd3293643094;
        test_addr[1697] = 471;
        test_data[1697] = 33'd1336088425;
        test_addr[1698] = 173;
        test_data[1698] = 33'd1456155483;
        test_addr[1699] = 854;
        test_data[1699] = 33'd2260897852;
        test_addr[1700] = 937;
        test_data[1700] = 33'd4794193628;
        test_addr[1701] = 316;
        test_data[1701] = 33'd3154340319;
        test_addr[1702] = 209;
        test_data[1702] = 33'd2185094724;
        test_addr[1703] = 661;
        test_data[1703] = 33'd5461807725;
        test_addr[1704] = 997;
        test_data[1704] = 33'd3981795757;
        test_addr[1705] = 788;
        test_data[1705] = 33'd3121816568;
        test_addr[1706] = 204;
        test_data[1706] = 33'd8243031507;
        test_addr[1707] = 773;
        test_data[1707] = 33'd1142927326;
        test_addr[1708] = 349;
        test_data[1708] = 33'd8215078497;
        test_addr[1709] = 47;
        test_data[1709] = 33'd1684233673;
        test_addr[1710] = 237;
        test_data[1710] = 33'd5346469526;
        test_addr[1711] = 853;
        test_data[1711] = 33'd3599534504;
        test_addr[1712] = 154;
        test_data[1712] = 33'd2265354610;
        test_addr[1713] = 839;
        test_data[1713] = 33'd709599084;
        test_addr[1714] = 573;
        test_data[1714] = 33'd5860187783;
        test_addr[1715] = 209;
        test_data[1715] = 33'd2185094724;
        test_addr[1716] = 793;
        test_data[1716] = 33'd1650429696;
        test_addr[1717] = 897;
        test_data[1717] = 33'd5079089413;
        test_addr[1718] = 720;
        test_data[1718] = 33'd713844621;
        test_addr[1719] = 329;
        test_data[1719] = 33'd3903899561;
        test_addr[1720] = 225;
        test_data[1720] = 33'd541535233;
        test_addr[1721] = 188;
        test_data[1721] = 33'd4083814239;
        test_addr[1722] = 777;
        test_data[1722] = 33'd1706937674;
        test_addr[1723] = 313;
        test_data[1723] = 33'd362309121;
        test_addr[1724] = 808;
        test_data[1724] = 33'd7789343176;
        test_addr[1725] = 705;
        test_data[1725] = 33'd5003835353;
        test_addr[1726] = 699;
        test_data[1726] = 33'd1968810960;
        test_addr[1727] = 871;
        test_data[1727] = 33'd6467390985;
        test_addr[1728] = 328;
        test_data[1728] = 33'd952282828;
        test_addr[1729] = 730;
        test_data[1729] = 33'd7126631442;
        test_addr[1730] = 199;
        test_data[1730] = 33'd1968015106;
        test_addr[1731] = 827;
        test_data[1731] = 33'd4136395276;
        test_addr[1732] = 157;
        test_data[1732] = 33'd1818871082;
        test_addr[1733] = 0;
        test_data[1733] = 33'd1940947903;
        test_addr[1734] = 199;
        test_data[1734] = 33'd1968015106;
        test_addr[1735] = 851;
        test_data[1735] = 33'd5067956094;
        test_addr[1736] = 769;
        test_data[1736] = 33'd3813893202;
        test_addr[1737] = 497;
        test_data[1737] = 33'd984535138;
        test_addr[1738] = 445;
        test_data[1738] = 33'd4845890257;
        test_addr[1739] = 207;
        test_data[1739] = 33'd843754471;
        test_addr[1740] = 905;
        test_data[1740] = 33'd2672417781;
        test_addr[1741] = 749;
        test_data[1741] = 33'd4915473940;
        test_addr[1742] = 446;
        test_data[1742] = 33'd1909467616;
        test_addr[1743] = 230;
        test_data[1743] = 33'd3123327297;
        test_addr[1744] = 765;
        test_data[1744] = 33'd1407724005;
        test_addr[1745] = 111;
        test_data[1745] = 33'd3462749259;
        test_addr[1746] = 615;
        test_data[1746] = 33'd2136755942;
        test_addr[1747] = 310;
        test_data[1747] = 33'd3692301779;
        test_addr[1748] = 857;
        test_data[1748] = 33'd1452427211;
        test_addr[1749] = 942;
        test_data[1749] = 33'd8486231303;
        test_addr[1750] = 67;
        test_data[1750] = 33'd3639768664;
        test_addr[1751] = 801;
        test_data[1751] = 33'd4743026103;
        test_addr[1752] = 268;
        test_data[1752] = 33'd6480595883;
        test_addr[1753] = 557;
        test_data[1753] = 33'd244671962;
        test_addr[1754] = 127;
        test_data[1754] = 33'd1731432911;
        test_addr[1755] = 674;
        test_data[1755] = 33'd2656360569;
        test_addr[1756] = 530;
        test_data[1756] = 33'd7311058765;
        test_addr[1757] = 265;
        test_data[1757] = 33'd3802763157;
        test_addr[1758] = 204;
        test_data[1758] = 33'd6587499895;
        test_addr[1759] = 732;
        test_data[1759] = 33'd3346690204;
        test_addr[1760] = 507;
        test_data[1760] = 33'd6724489436;
        test_addr[1761] = 966;
        test_data[1761] = 33'd1835137690;
        test_addr[1762] = 785;
        test_data[1762] = 33'd1401173062;
        test_addr[1763] = 34;
        test_data[1763] = 33'd2988630753;
        test_addr[1764] = 909;
        test_data[1764] = 33'd3935995031;
        test_addr[1765] = 610;
        test_data[1765] = 33'd6270289556;
        test_addr[1766] = 938;
        test_data[1766] = 33'd6583595422;
        test_addr[1767] = 229;
        test_data[1767] = 33'd920626449;
        test_addr[1768] = 102;
        test_data[1768] = 33'd1124317209;
        test_addr[1769] = 121;
        test_data[1769] = 33'd157354656;
        test_addr[1770] = 134;
        test_data[1770] = 33'd2206256073;
        test_addr[1771] = 80;
        test_data[1771] = 33'd818068638;
        test_addr[1772] = 952;
        test_data[1772] = 33'd702855526;
        test_addr[1773] = 469;
        test_data[1773] = 33'd3211600796;
        test_addr[1774] = 189;
        test_data[1774] = 33'd3994613051;
        test_addr[1775] = 136;
        test_data[1775] = 33'd3019476229;
        test_addr[1776] = 226;
        test_data[1776] = 33'd5561350609;
        test_addr[1777] = 215;
        test_data[1777] = 33'd8030626571;
        test_addr[1778] = 333;
        test_data[1778] = 33'd5125370450;
        test_addr[1779] = 31;
        test_data[1779] = 33'd1855015640;
        test_addr[1780] = 616;
        test_data[1780] = 33'd4761171635;
        test_addr[1781] = 512;
        test_data[1781] = 33'd112430786;
        test_addr[1782] = 10;
        test_data[1782] = 33'd3594809116;
        test_addr[1783] = 410;
        test_data[1783] = 33'd3405405453;
        test_addr[1784] = 793;
        test_data[1784] = 33'd1650429696;
        test_addr[1785] = 818;
        test_data[1785] = 33'd3872489273;
        test_addr[1786] = 773;
        test_data[1786] = 33'd1142927326;
        test_addr[1787] = 716;
        test_data[1787] = 33'd1341092090;
        test_addr[1788] = 648;
        test_data[1788] = 33'd5231450239;
        test_addr[1789] = 909;
        test_data[1789] = 33'd7491916262;
        test_addr[1790] = 363;
        test_data[1790] = 33'd7293023377;
        test_addr[1791] = 631;
        test_data[1791] = 33'd6811379858;
        test_addr[1792] = 566;
        test_data[1792] = 33'd7888820663;
        test_addr[1793] = 884;
        test_data[1793] = 33'd1323552558;
        test_addr[1794] = 389;
        test_data[1794] = 33'd2549642068;
        test_addr[1795] = 544;
        test_data[1795] = 33'd7450513492;
        test_addr[1796] = 212;
        test_data[1796] = 33'd1617687132;
        test_addr[1797] = 485;
        test_data[1797] = 33'd1200863765;
        test_addr[1798] = 571;
        test_data[1798] = 33'd3849053210;
        test_addr[1799] = 61;
        test_data[1799] = 33'd5588221606;
        test_addr[1800] = 865;
        test_data[1800] = 33'd6797875861;
        test_addr[1801] = 662;
        test_data[1801] = 33'd2183779360;
        test_addr[1802] = 535;
        test_data[1802] = 33'd1384824159;
        test_addr[1803] = 465;
        test_data[1803] = 33'd896820312;
        test_addr[1804] = 219;
        test_data[1804] = 33'd308900539;
        test_addr[1805] = 943;
        test_data[1805] = 33'd6070364149;
        test_addr[1806] = 858;
        test_data[1806] = 33'd1025625720;
        test_addr[1807] = 779;
        test_data[1807] = 33'd2260017456;
        test_addr[1808] = 825;
        test_data[1808] = 33'd1248929761;
        test_addr[1809] = 530;
        test_data[1809] = 33'd3016091469;
        test_addr[1810] = 717;
        test_data[1810] = 33'd2102291868;
        test_addr[1811] = 781;
        test_data[1811] = 33'd2061765198;
        test_addr[1812] = 510;
        test_data[1812] = 33'd363583401;
        test_addr[1813] = 314;
        test_data[1813] = 33'd5003828054;
        test_addr[1814] = 876;
        test_data[1814] = 33'd2922270056;
        test_addr[1815] = 881;
        test_data[1815] = 33'd554101517;
        test_addr[1816] = 393;
        test_data[1816] = 33'd7355044714;
        test_addr[1817] = 588;
        test_data[1817] = 33'd4041263385;
        test_addr[1818] = 604;
        test_data[1818] = 33'd70723367;
        test_addr[1819] = 315;
        test_data[1819] = 33'd3577492034;
        test_addr[1820] = 387;
        test_data[1820] = 33'd984172897;
        test_addr[1821] = 509;
        test_data[1821] = 33'd3789326765;
        test_addr[1822] = 366;
        test_data[1822] = 33'd648433376;
        test_addr[1823] = 789;
        test_data[1823] = 33'd2899379877;
        test_addr[1824] = 378;
        test_data[1824] = 33'd7264099384;
        test_addr[1825] = 998;
        test_data[1825] = 33'd3897224364;
        test_addr[1826] = 453;
        test_data[1826] = 33'd6856674125;
        test_addr[1827] = 480;
        test_data[1827] = 33'd648309832;
        test_addr[1828] = 656;
        test_data[1828] = 33'd2637048261;
        test_addr[1829] = 220;
        test_data[1829] = 33'd1136133958;
        test_addr[1830] = 982;
        test_data[1830] = 33'd7324085184;
        test_addr[1831] = 23;
        test_data[1831] = 33'd1087399442;
        test_addr[1832] = 556;
        test_data[1832] = 33'd2030797940;
        test_addr[1833] = 148;
        test_data[1833] = 33'd1899923406;
        test_addr[1834] = 915;
        test_data[1834] = 33'd1268898235;
        test_addr[1835] = 654;
        test_data[1835] = 33'd1773452330;
        test_addr[1836] = 932;
        test_data[1836] = 33'd8570095673;
        test_addr[1837] = 720;
        test_data[1837] = 33'd5531868359;
        test_addr[1838] = 66;
        test_data[1838] = 33'd5815587083;
        test_addr[1839] = 564;
        test_data[1839] = 33'd2953020563;
        test_addr[1840] = 583;
        test_data[1840] = 33'd1888552959;
        test_addr[1841] = 918;
        test_data[1841] = 33'd2681524291;
        test_addr[1842] = 114;
        test_data[1842] = 33'd4780989762;
        test_addr[1843] = 91;
        test_data[1843] = 33'd8168171827;
        test_addr[1844] = 249;
        test_data[1844] = 33'd8289272830;
        test_addr[1845] = 329;
        test_data[1845] = 33'd6747962430;
        test_addr[1846] = 696;
        test_data[1846] = 33'd2694337344;
        test_addr[1847] = 318;
        test_data[1847] = 33'd1218864492;
        test_addr[1848] = 361;
        test_data[1848] = 33'd3444719037;
        test_addr[1849] = 605;
        test_data[1849] = 33'd1980249529;
        test_addr[1850] = 502;
        test_data[1850] = 33'd5752738270;
        test_addr[1851] = 148;
        test_data[1851] = 33'd4419846177;
        test_addr[1852] = 896;
        test_data[1852] = 33'd3625741568;
        test_addr[1853] = 824;
        test_data[1853] = 33'd311419234;
        test_addr[1854] = 642;
        test_data[1854] = 33'd4370365240;
        test_addr[1855] = 540;
        test_data[1855] = 33'd432267239;
        test_addr[1856] = 901;
        test_data[1856] = 33'd3791968021;
        test_addr[1857] = 595;
        test_data[1857] = 33'd8129462238;
        test_addr[1858] = 40;
        test_data[1858] = 33'd2224301287;
        test_addr[1859] = 660;
        test_data[1859] = 33'd1826723096;
        test_addr[1860] = 132;
        test_data[1860] = 33'd3529417599;
        test_addr[1861] = 75;
        test_data[1861] = 33'd2274537304;
        test_addr[1862] = 471;
        test_data[1862] = 33'd4890107594;
        test_addr[1863] = 579;
        test_data[1863] = 33'd2718604588;
        test_addr[1864] = 29;
        test_data[1864] = 33'd131073219;
        test_addr[1865] = 395;
        test_data[1865] = 33'd1292390397;
        test_addr[1866] = 1023;
        test_data[1866] = 33'd4626912356;
        test_addr[1867] = 54;
        test_data[1867] = 33'd559000320;
        test_addr[1868] = 16;
        test_data[1868] = 33'd6528664110;
        test_addr[1869] = 260;
        test_data[1869] = 33'd5812919125;
        test_addr[1870] = 87;
        test_data[1870] = 33'd3922461656;
        test_addr[1871] = 979;
        test_data[1871] = 33'd4346784549;
        test_addr[1872] = 186;
        test_data[1872] = 33'd1670278583;
        test_addr[1873] = 163;
        test_data[1873] = 33'd6517198163;
        test_addr[1874] = 868;
        test_data[1874] = 33'd2528507951;
        test_addr[1875] = 562;
        test_data[1875] = 33'd4108954016;
        test_addr[1876] = 240;
        test_data[1876] = 33'd3107113144;
        test_addr[1877] = 400;
        test_data[1877] = 33'd545504374;
        test_addr[1878] = 678;
        test_data[1878] = 33'd2022273082;
        test_addr[1879] = 622;
        test_data[1879] = 33'd3351421963;
        test_addr[1880] = 337;
        test_data[1880] = 33'd6921767378;
        test_addr[1881] = 393;
        test_data[1881] = 33'd5308472386;
        test_addr[1882] = 226;
        test_data[1882] = 33'd6832647763;
        test_addr[1883] = 554;
        test_data[1883] = 33'd2207183766;
        test_addr[1884] = 832;
        test_data[1884] = 33'd351971474;
        test_addr[1885] = 818;
        test_data[1885] = 33'd4997375713;
        test_addr[1886] = 283;
        test_data[1886] = 33'd581010001;
        test_addr[1887] = 683;
        test_data[1887] = 33'd8289489171;
        test_addr[1888] = 12;
        test_data[1888] = 33'd4028186270;
        test_addr[1889] = 754;
        test_data[1889] = 33'd1231791903;
        test_addr[1890] = 292;
        test_data[1890] = 33'd7114363558;
        test_addr[1891] = 342;
        test_data[1891] = 33'd6109849748;
        test_addr[1892] = 137;
        test_data[1892] = 33'd8101690043;
        test_addr[1893] = 764;
        test_data[1893] = 33'd82671605;
        test_addr[1894] = 851;
        test_data[1894] = 33'd6392259657;
        test_addr[1895] = 250;
        test_data[1895] = 33'd673588786;
        test_addr[1896] = 815;
        test_data[1896] = 33'd1640602374;
        test_addr[1897] = 322;
        test_data[1897] = 33'd3243207308;
        test_addr[1898] = 796;
        test_data[1898] = 33'd4142487238;
        test_addr[1899] = 246;
        test_data[1899] = 33'd1635138116;
        test_addr[1900] = 745;
        test_data[1900] = 33'd469000044;
        test_addr[1901] = 258;
        test_data[1901] = 33'd2974304192;
        test_addr[1902] = 848;
        test_data[1902] = 33'd6679614770;
        test_addr[1903] = 924;
        test_data[1903] = 33'd2714813433;
        test_addr[1904] = 834;
        test_data[1904] = 33'd1152692795;
        test_addr[1905] = 802;
        test_data[1905] = 33'd8239738986;
        test_addr[1906] = 403;
        test_data[1906] = 33'd2351946442;
        test_addr[1907] = 406;
        test_data[1907] = 33'd1667658830;
        test_addr[1908] = 541;
        test_data[1908] = 33'd4208840303;
        test_addr[1909] = 727;
        test_data[1909] = 33'd8355975047;
        test_addr[1910] = 394;
        test_data[1910] = 33'd1231576489;
        test_addr[1911] = 759;
        test_data[1911] = 33'd6491847183;
        test_addr[1912] = 271;
        test_data[1912] = 33'd4939598316;
        test_addr[1913] = 92;
        test_data[1913] = 33'd1230523681;
        test_addr[1914] = 546;
        test_data[1914] = 33'd4850769435;
        test_addr[1915] = 110;
        test_data[1915] = 33'd916244885;
        test_addr[1916] = 674;
        test_data[1916] = 33'd2656360569;
        test_addr[1917] = 471;
        test_data[1917] = 33'd595140298;
        test_addr[1918] = 835;
        test_data[1918] = 33'd6424899992;
        test_addr[1919] = 680;
        test_data[1919] = 33'd5179049369;
        test_addr[1920] = 27;
        test_data[1920] = 33'd5165071535;
        test_addr[1921] = 500;
        test_data[1921] = 33'd7159532380;
        test_addr[1922] = 194;
        test_data[1922] = 33'd2912051046;
        test_addr[1923] = 51;
        test_data[1923] = 33'd1434736929;
        test_addr[1924] = 158;
        test_data[1924] = 33'd217812934;
        test_addr[1925] = 63;
        test_data[1925] = 33'd2633027552;
        test_addr[1926] = 157;
        test_data[1926] = 33'd6812015773;
        test_addr[1927] = 935;
        test_data[1927] = 33'd8153228866;
        test_addr[1928] = 305;
        test_data[1928] = 33'd1101688979;
        test_addr[1929] = 498;
        test_data[1929] = 33'd3649231511;
        test_addr[1930] = 222;
        test_data[1930] = 33'd8079629613;
        test_addr[1931] = 848;
        test_data[1931] = 33'd2384647474;
        test_addr[1932] = 350;
        test_data[1932] = 33'd3976893991;
        test_addr[1933] = 404;
        test_data[1933] = 33'd214098716;
        test_addr[1934] = 249;
        test_data[1934] = 33'd3994305534;
        test_addr[1935] = 845;
        test_data[1935] = 33'd1963746399;
        test_addr[1936] = 266;
        test_data[1936] = 33'd4693562488;
        test_addr[1937] = 987;
        test_data[1937] = 33'd5656762299;
        test_addr[1938] = 488;
        test_data[1938] = 33'd5134648100;
        test_addr[1939] = 203;
        test_data[1939] = 33'd4132021586;
        test_addr[1940] = 1016;
        test_data[1940] = 33'd6221751970;
        test_addr[1941] = 927;
        test_data[1941] = 33'd1927721038;
        test_addr[1942] = 417;
        test_data[1942] = 33'd2268883569;
        test_addr[1943] = 155;
        test_data[1943] = 33'd1302683176;
        test_addr[1944] = 958;
        test_data[1944] = 33'd3257284543;
        test_addr[1945] = 904;
        test_data[1945] = 33'd580095324;
        test_addr[1946] = 790;
        test_data[1946] = 33'd7343677487;
        test_addr[1947] = 70;
        test_data[1947] = 33'd1368704711;
        test_addr[1948] = 133;
        test_data[1948] = 33'd4790786856;
        test_addr[1949] = 617;
        test_data[1949] = 33'd2620405328;
        test_addr[1950] = 239;
        test_data[1950] = 33'd1377847727;
        test_addr[1951] = 260;
        test_data[1951] = 33'd1517951829;
        test_addr[1952] = 945;
        test_data[1952] = 33'd4667001816;
        test_addr[1953] = 255;
        test_data[1953] = 33'd1916824779;
        test_addr[1954] = 857;
        test_data[1954] = 33'd1452427211;
        test_addr[1955] = 908;
        test_data[1955] = 33'd5999821660;
        test_addr[1956] = 823;
        test_data[1956] = 33'd1932951958;
        test_addr[1957] = 46;
        test_data[1957] = 33'd4095908597;
        test_addr[1958] = 807;
        test_data[1958] = 33'd4145466213;
        test_addr[1959] = 1022;
        test_data[1959] = 33'd7545942847;
        test_addr[1960] = 1005;
        test_data[1960] = 33'd1098300837;
        test_addr[1961] = 390;
        test_data[1961] = 33'd909123417;
        test_addr[1962] = 501;
        test_data[1962] = 33'd3623861933;
        test_addr[1963] = 696;
        test_data[1963] = 33'd2694337344;
        test_addr[1964] = 728;
        test_data[1964] = 33'd806584098;
        test_addr[1965] = 590;
        test_data[1965] = 33'd254542356;
        test_addr[1966] = 239;
        test_data[1966] = 33'd1377847727;
        test_addr[1967] = 582;
        test_data[1967] = 33'd5822564396;
        test_addr[1968] = 792;
        test_data[1968] = 33'd4103913134;
        test_addr[1969] = 339;
        test_data[1969] = 33'd232710529;
        test_addr[1970] = 931;
        test_data[1970] = 33'd2803979244;
        test_addr[1971] = 518;
        test_data[1971] = 33'd6801143411;
        test_addr[1972] = 442;
        test_data[1972] = 33'd7816694134;
        test_addr[1973] = 925;
        test_data[1973] = 33'd7991977669;
        test_addr[1974] = 857;
        test_data[1974] = 33'd5615571775;
        test_addr[1975] = 60;
        test_data[1975] = 33'd7989653969;
        test_addr[1976] = 50;
        test_data[1976] = 33'd1433122672;
        test_addr[1977] = 578;
        test_data[1977] = 33'd1262376951;
        test_addr[1978] = 93;
        test_data[1978] = 33'd5811643138;
        test_addr[1979] = 927;
        test_data[1979] = 33'd7176618952;
        test_addr[1980] = 980;
        test_data[1980] = 33'd3594942886;
        test_addr[1981] = 106;
        test_data[1981] = 33'd898134430;
        test_addr[1982] = 780;
        test_data[1982] = 33'd404411201;
        test_addr[1983] = 852;
        test_data[1983] = 33'd4803826115;
        test_addr[1984] = 854;
        test_data[1984] = 33'd2260897852;
        test_addr[1985] = 491;
        test_data[1985] = 33'd8064909174;
        test_addr[1986] = 651;
        test_data[1986] = 33'd1359098933;
        test_addr[1987] = 840;
        test_data[1987] = 33'd788849187;
        test_addr[1988] = 699;
        test_data[1988] = 33'd1968810960;
        test_addr[1989] = 387;
        test_data[1989] = 33'd7359743551;
        test_addr[1990] = 381;
        test_data[1990] = 33'd1838811245;
        test_addr[1991] = 1021;
        test_data[1991] = 33'd1393906874;
        test_addr[1992] = 354;
        test_data[1992] = 33'd2820300650;
        test_addr[1993] = 952;
        test_data[1993] = 33'd8368156359;
        test_addr[1994] = 96;
        test_data[1994] = 33'd3127743323;
        test_addr[1995] = 690;
        test_data[1995] = 33'd4095690594;
        test_addr[1996] = 437;
        test_data[1996] = 33'd3188866646;
        test_addr[1997] = 285;
        test_data[1997] = 33'd5861757806;
        test_addr[1998] = 160;
        test_data[1998] = 33'd772555075;
        test_addr[1999] = 677;
        test_data[1999] = 33'd7280132683;
        test_addr[2000] = 52;
        test_data[2000] = 33'd7889071808;
        test_addr[2001] = 769;
        test_data[2001] = 33'd3813893202;
        test_addr[2002] = 595;
        test_data[2002] = 33'd4560385130;
        test_addr[2003] = 29;
        test_data[2003] = 33'd4555161106;
        test_addr[2004] = 467;
        test_data[2004] = 33'd2928862965;
        test_addr[2005] = 454;
        test_data[2005] = 33'd3130965914;
        test_addr[2006] = 520;
        test_data[2006] = 33'd4312066109;
        test_addr[2007] = 992;
        test_data[2007] = 33'd3283916326;
        test_addr[2008] = 969;
        test_data[2008] = 33'd5927331253;
        test_addr[2009] = 707;
        test_data[2009] = 33'd866118162;
        test_addr[2010] = 22;
        test_data[2010] = 33'd9397193;
        test_addr[2011] = 424;
        test_data[2011] = 33'd710281784;
        test_addr[2012] = 404;
        test_data[2012] = 33'd214098716;
        test_addr[2013] = 730;
        test_data[2013] = 33'd8508652960;
        test_addr[2014] = 300;
        test_data[2014] = 33'd4668844694;
        test_addr[2015] = 935;
        test_data[2015] = 33'd3858261570;
        test_addr[2016] = 221;
        test_data[2016] = 33'd720358563;
        test_addr[2017] = 884;
        test_data[2017] = 33'd1323552558;
        test_addr[2018] = 590;
        test_data[2018] = 33'd254542356;
        test_addr[2019] = 942;
        test_data[2019] = 33'd6144661171;
        test_addr[2020] = 718;
        test_data[2020] = 33'd2587264415;
        test_addr[2021] = 1015;
        test_data[2021] = 33'd2062647632;
        test_addr[2022] = 754;
        test_data[2022] = 33'd1231791903;
        test_addr[2023] = 817;
        test_data[2023] = 33'd5089817717;
        test_addr[2024] = 291;
        test_data[2024] = 33'd4584240249;
        test_addr[2025] = 1014;
        test_data[2025] = 33'd7831124607;
        test_addr[2026] = 377;
        test_data[2026] = 33'd2370864657;
        test_addr[2027] = 138;
        test_data[2027] = 33'd2910298998;
        test_addr[2028] = 48;
        test_data[2028] = 33'd3748276960;
        test_addr[2029] = 1020;
        test_data[2029] = 33'd1993492834;
        test_addr[2030] = 272;
        test_data[2030] = 33'd478200901;
        test_addr[2031] = 882;
        test_data[2031] = 33'd4205936978;
        test_addr[2032] = 92;
        test_data[2032] = 33'd1230523681;
        test_addr[2033] = 42;
        test_data[2033] = 33'd3652372969;
        test_addr[2034] = 791;
        test_data[2034] = 33'd1738721985;
        test_addr[2035] = 58;
        test_data[2035] = 33'd4758603810;
        test_addr[2036] = 509;
        test_data[2036] = 33'd7426736617;
        test_addr[2037] = 522;
        test_data[2037] = 33'd5800478481;
        test_addr[2038] = 978;
        test_data[2038] = 33'd1609416996;
        test_addr[2039] = 722;
        test_data[2039] = 33'd5522443214;
        test_addr[2040] = 973;
        test_data[2040] = 33'd986805218;
        test_addr[2041] = 811;
        test_data[2041] = 33'd712960676;
        test_addr[2042] = 154;
        test_data[2042] = 33'd2265354610;
        test_addr[2043] = 705;
        test_data[2043] = 33'd7380510414;
        test_addr[2044] = 39;
        test_data[2044] = 33'd3634135297;
        test_addr[2045] = 347;
        test_data[2045] = 33'd3874808649;
        test_addr[2046] = 1005;
        test_data[2046] = 33'd1098300837;
        test_addr[2047] = 603;
        test_data[2047] = 33'd2447831809;
        test_addr[2048] = 455;
        test_data[2048] = 33'd2867352729;
        test_addr[2049] = 573;
        test_data[2049] = 33'd1565220487;
        test_addr[2050] = 617;
        test_data[2050] = 33'd5178902897;
        test_addr[2051] = 680;
        test_data[2051] = 33'd884082073;
        test_addr[2052] = 244;
        test_data[2052] = 33'd656960195;
        test_addr[2053] = 273;
        test_data[2053] = 33'd56693191;
        test_addr[2054] = 337;
        test_data[2054] = 33'd2626800082;
        test_addr[2055] = 692;
        test_data[2055] = 33'd366443818;
        test_addr[2056] = 217;
        test_data[2056] = 33'd8199352024;
        test_addr[2057] = 336;
        test_data[2057] = 33'd2382706043;
        test_addr[2058] = 827;
        test_data[2058] = 33'd4136395276;
        test_addr[2059] = 369;
        test_data[2059] = 33'd7057348042;
        test_addr[2060] = 627;
        test_data[2060] = 33'd6173483377;
        test_addr[2061] = 340;
        test_data[2061] = 33'd3309872861;
        test_addr[2062] = 365;
        test_data[2062] = 33'd369210451;
        test_addr[2063] = 320;
        test_data[2063] = 33'd7870305742;
        test_addr[2064] = 128;
        test_data[2064] = 33'd7968480493;
        test_addr[2065] = 887;
        test_data[2065] = 33'd6675657320;
        test_addr[2066] = 207;
        test_data[2066] = 33'd5087803885;
        test_addr[2067] = 20;
        test_data[2067] = 33'd4222788375;
        test_addr[2068] = 983;
        test_data[2068] = 33'd509354105;
        test_addr[2069] = 712;
        test_data[2069] = 33'd1104352139;
        test_addr[2070] = 585;
        test_data[2070] = 33'd3586969900;
        test_addr[2071] = 784;
        test_data[2071] = 33'd4161914853;
        test_addr[2072] = 695;
        test_data[2072] = 33'd2186911345;
        test_addr[2073] = 294;
        test_data[2073] = 33'd228860212;
        test_addr[2074] = 328;
        test_data[2074] = 33'd952282828;
        test_addr[2075] = 837;
        test_data[2075] = 33'd2747873873;
        test_addr[2076] = 962;
        test_data[2076] = 33'd3905065194;
        test_addr[2077] = 584;
        test_data[2077] = 33'd3681182924;
        test_addr[2078] = 865;
        test_data[2078] = 33'd2502908565;
        test_addr[2079] = 705;
        test_data[2079] = 33'd3085543118;
        test_addr[2080] = 233;
        test_data[2080] = 33'd1289878889;
        test_addr[2081] = 857;
        test_data[2081] = 33'd1320604479;
        test_addr[2082] = 327;
        test_data[2082] = 33'd6307703250;
        test_addr[2083] = 740;
        test_data[2083] = 33'd1790213294;
        test_addr[2084] = 1017;
        test_data[2084] = 33'd7943649734;
        test_addr[2085] = 453;
        test_data[2085] = 33'd2561706829;
        test_addr[2086] = 736;
        test_data[2086] = 33'd1931613996;
        test_addr[2087] = 315;
        test_data[2087] = 33'd3577492034;
        test_addr[2088] = 585;
        test_data[2088] = 33'd3586969900;
        test_addr[2089] = 220;
        test_data[2089] = 33'd1136133958;
        test_addr[2090] = 253;
        test_data[2090] = 33'd2796634323;
        test_addr[2091] = 517;
        test_data[2091] = 33'd385111081;
        test_addr[2092] = 659;
        test_data[2092] = 33'd2764015169;
        test_addr[2093] = 849;
        test_data[2093] = 33'd7615520888;
        test_addr[2094] = 64;
        test_data[2094] = 33'd3038722049;
        test_addr[2095] = 954;
        test_data[2095] = 33'd1594670622;
        test_addr[2096] = 172;
        test_data[2096] = 33'd1555194164;
        test_addr[2097] = 541;
        test_data[2097] = 33'd4208840303;
        test_addr[2098] = 384;
        test_data[2098] = 33'd4961229841;
        test_addr[2099] = 628;
        test_data[2099] = 33'd8197680955;
        test_addr[2100] = 156;
        test_data[2100] = 33'd3852022963;
        test_addr[2101] = 694;
        test_data[2101] = 33'd240080374;
        test_addr[2102] = 591;
        test_data[2102] = 33'd7701701295;
        test_addr[2103] = 869;
        test_data[2103] = 33'd2336492666;
        test_addr[2104] = 199;
        test_data[2104] = 33'd1968015106;
        test_addr[2105] = 347;
        test_data[2105] = 33'd3874808649;
        test_addr[2106] = 375;
        test_data[2106] = 33'd1408822660;
        test_addr[2107] = 890;
        test_data[2107] = 33'd2018427355;
        test_addr[2108] = 716;
        test_data[2108] = 33'd7398385203;
        test_addr[2109] = 1022;
        test_data[2109] = 33'd3250975551;
        test_addr[2110] = 717;
        test_data[2110] = 33'd2102291868;
        test_addr[2111] = 109;
        test_data[2111] = 33'd2394762171;
        test_addr[2112] = 942;
        test_data[2112] = 33'd6428708952;
        test_addr[2113] = 601;
        test_data[2113] = 33'd2919076942;
        test_addr[2114] = 798;
        test_data[2114] = 33'd4195757002;
        test_addr[2115] = 310;
        test_data[2115] = 33'd3692301779;
        test_addr[2116] = 371;
        test_data[2116] = 33'd941454407;
        test_addr[2117] = 25;
        test_data[2117] = 33'd2605255280;
        test_addr[2118] = 2;
        test_data[2118] = 33'd3771999802;
        test_addr[2119] = 925;
        test_data[2119] = 33'd3697010373;
        test_addr[2120] = 774;
        test_data[2120] = 33'd197646308;
        test_addr[2121] = 300;
        test_data[2121] = 33'd6420272191;
        test_addr[2122] = 719;
        test_data[2122] = 33'd3780764175;
        test_addr[2123] = 749;
        test_data[2123] = 33'd5282403148;
        test_addr[2124] = 405;
        test_data[2124] = 33'd516109638;
        test_addr[2125] = 913;
        test_data[2125] = 33'd2312966920;
        test_addr[2126] = 888;
        test_data[2126] = 33'd1386718648;
        test_addr[2127] = 398;
        test_data[2127] = 33'd1175204693;
        test_addr[2128] = 989;
        test_data[2128] = 33'd2812472571;
        test_addr[2129] = 741;
        test_data[2129] = 33'd3239258243;
        test_addr[2130] = 608;
        test_data[2130] = 33'd3381739994;
        test_addr[2131] = 528;
        test_data[2131] = 33'd3121538625;
        test_addr[2132] = 101;
        test_data[2132] = 33'd5304358273;
        test_addr[2133] = 408;
        test_data[2133] = 33'd1130836166;
        test_addr[2134] = 312;
        test_data[2134] = 33'd7006609782;
        test_addr[2135] = 717;
        test_data[2135] = 33'd8176267513;
        test_addr[2136] = 534;
        test_data[2136] = 33'd2464887914;
        test_addr[2137] = 468;
        test_data[2137] = 33'd49837857;
        test_addr[2138] = 730;
        test_data[2138] = 33'd4658048373;
        test_addr[2139] = 594;
        test_data[2139] = 33'd7230905202;
        test_addr[2140] = 866;
        test_data[2140] = 33'd3574629408;
        test_addr[2141] = 477;
        test_data[2141] = 33'd5379841529;
        test_addr[2142] = 733;
        test_data[2142] = 33'd3710281497;
        test_addr[2143] = 625;
        test_data[2143] = 33'd4896798263;
        test_addr[2144] = 947;
        test_data[2144] = 33'd4717100386;
        test_addr[2145] = 482;
        test_data[2145] = 33'd7100257272;
        test_addr[2146] = 332;
        test_data[2146] = 33'd2406902933;
        test_addr[2147] = 699;
        test_data[2147] = 33'd1968810960;
        test_addr[2148] = 520;
        test_data[2148] = 33'd8308061304;
        test_addr[2149] = 539;
        test_data[2149] = 33'd6925771774;
        test_addr[2150] = 201;
        test_data[2150] = 33'd29735866;
        test_addr[2151] = 624;
        test_data[2151] = 33'd3776573770;
        test_addr[2152] = 768;
        test_data[2152] = 33'd3795726059;
        test_addr[2153] = 679;
        test_data[2153] = 33'd8170110300;
        test_addr[2154] = 300;
        test_data[2154] = 33'd4827492055;
        test_addr[2155] = 323;
        test_data[2155] = 33'd1032448390;
        test_addr[2156] = 116;
        test_data[2156] = 33'd5215594401;
        test_addr[2157] = 690;
        test_data[2157] = 33'd4095690594;
        test_addr[2158] = 718;
        test_data[2158] = 33'd2587264415;
        test_addr[2159] = 331;
        test_data[2159] = 33'd3237563871;
        test_addr[2160] = 203;
        test_data[2160] = 33'd6972267689;
        test_addr[2161] = 52;
        test_data[2161] = 33'd3594104512;
        test_addr[2162] = 56;
        test_data[2162] = 33'd3847507083;
        test_addr[2163] = 1013;
        test_data[2163] = 33'd519919884;
        test_addr[2164] = 539;
        test_data[2164] = 33'd8106797100;
        test_addr[2165] = 800;
        test_data[2165] = 33'd2470310901;
        test_addr[2166] = 475;
        test_data[2166] = 33'd7309859880;
        test_addr[2167] = 55;
        test_data[2167] = 33'd4289280957;
        test_addr[2168] = 970;
        test_data[2168] = 33'd5043913511;
        test_addr[2169] = 861;
        test_data[2169] = 33'd7615436071;
        test_addr[2170] = 177;
        test_data[2170] = 33'd2198187797;
        test_addr[2171] = 202;
        test_data[2171] = 33'd1530277351;
        test_addr[2172] = 56;
        test_data[2172] = 33'd3847507083;
        test_addr[2173] = 705;
        test_data[2173] = 33'd5771752300;
        test_addr[2174] = 951;
        test_data[2174] = 33'd4806602225;
        test_addr[2175] = 367;
        test_data[2175] = 33'd5856786932;
        test_addr[2176] = 973;
        test_data[2176] = 33'd986805218;
        test_addr[2177] = 504;
        test_data[2177] = 33'd2373341895;
        test_addr[2178] = 658;
        test_data[2178] = 33'd7197369872;
        test_addr[2179] = 616;
        test_data[2179] = 33'd466204339;
        test_addr[2180] = 651;
        test_data[2180] = 33'd6505852862;
        test_addr[2181] = 79;
        test_data[2181] = 33'd8059009511;
        test_addr[2182] = 940;
        test_data[2182] = 33'd2857151879;
        test_addr[2183] = 534;
        test_data[2183] = 33'd2464887914;
        test_addr[2184] = 597;
        test_data[2184] = 33'd7442783782;
        test_addr[2185] = 484;
        test_data[2185] = 33'd953158137;
        test_addr[2186] = 476;
        test_data[2186] = 33'd8143470933;
        test_addr[2187] = 201;
        test_data[2187] = 33'd29735866;
        test_addr[2188] = 335;
        test_data[2188] = 33'd2081762056;
        test_addr[2189] = 515;
        test_data[2189] = 33'd1989592525;
        test_addr[2190] = 441;
        test_data[2190] = 33'd1603229292;
        test_addr[2191] = 29;
        test_data[2191] = 33'd260193810;
        test_addr[2192] = 957;
        test_data[2192] = 33'd7165897081;
        test_addr[2193] = 977;
        test_data[2193] = 33'd1687923687;
        test_addr[2194] = 651;
        test_data[2194] = 33'd2210885566;
        test_addr[2195] = 371;
        test_data[2195] = 33'd941454407;
        test_addr[2196] = 345;
        test_data[2196] = 33'd2662284645;
        test_addr[2197] = 873;
        test_data[2197] = 33'd722926779;
        test_addr[2198] = 900;
        test_data[2198] = 33'd3715729542;
        test_addr[2199] = 920;
        test_data[2199] = 33'd7398686110;
        test_addr[2200] = 252;
        test_data[2200] = 33'd1173487842;
        test_addr[2201] = 543;
        test_data[2201] = 33'd3369326361;
        test_addr[2202] = 101;
        test_data[2202] = 33'd7567399468;
        test_addr[2203] = 808;
        test_data[2203] = 33'd3494375880;
        test_addr[2204] = 533;
        test_data[2204] = 33'd3809017245;
        test_addr[2205] = 592;
        test_data[2205] = 33'd938793682;
        test_addr[2206] = 293;
        test_data[2206] = 33'd5954165169;
        test_addr[2207] = 160;
        test_data[2207] = 33'd772555075;
        test_addr[2208] = 337;
        test_data[2208] = 33'd2626800082;
        test_addr[2209] = 796;
        test_data[2209] = 33'd4142487238;
        test_addr[2210] = 661;
        test_data[2210] = 33'd1166840429;
        test_addr[2211] = 522;
        test_data[2211] = 33'd7741019135;
        test_addr[2212] = 959;
        test_data[2212] = 33'd910132403;
        test_addr[2213] = 558;
        test_data[2213] = 33'd3650811963;
        test_addr[2214] = 458;
        test_data[2214] = 33'd3114864730;
        test_addr[2215] = 528;
        test_data[2215] = 33'd7956758240;
        test_addr[2216] = 473;
        test_data[2216] = 33'd8416888412;
        test_addr[2217] = 834;
        test_data[2217] = 33'd7399694961;
        test_addr[2218] = 270;
        test_data[2218] = 33'd6517380875;
        test_addr[2219] = 247;
        test_data[2219] = 33'd4009011063;
        test_addr[2220] = 895;
        test_data[2220] = 33'd2337862672;
        test_addr[2221] = 280;
        test_data[2221] = 33'd1449766228;
        test_addr[2222] = 427;
        test_data[2222] = 33'd3998550133;
        test_addr[2223] = 132;
        test_data[2223] = 33'd3529417599;
        test_addr[2224] = 746;
        test_data[2224] = 33'd2332255621;
        test_addr[2225] = 462;
        test_data[2225] = 33'd3869809521;
        test_addr[2226] = 469;
        test_data[2226] = 33'd3211600796;
        test_addr[2227] = 852;
        test_data[2227] = 33'd5353757691;
        test_addr[2228] = 399;
        test_data[2228] = 33'd4989071036;
        test_addr[2229] = 1018;
        test_data[2229] = 33'd2731182889;
        test_addr[2230] = 631;
        test_data[2230] = 33'd6165169560;
        test_addr[2231] = 322;
        test_data[2231] = 33'd3243207308;
        test_addr[2232] = 313;
        test_data[2232] = 33'd6400604876;
        test_addr[2233] = 523;
        test_data[2233] = 33'd577685601;
        test_addr[2234] = 377;
        test_data[2234] = 33'd2370864657;
        test_addr[2235] = 270;
        test_data[2235] = 33'd2222413579;
        test_addr[2236] = 433;
        test_data[2236] = 33'd4722848486;
        test_addr[2237] = 562;
        test_data[2237] = 33'd4874056998;
        test_addr[2238] = 876;
        test_data[2238] = 33'd2922270056;
        test_addr[2239] = 395;
        test_data[2239] = 33'd7737093911;
        test_addr[2240] = 429;
        test_data[2240] = 33'd2701848083;
        test_addr[2241] = 788;
        test_data[2241] = 33'd3121816568;
        test_addr[2242] = 834;
        test_data[2242] = 33'd3104727665;
        test_addr[2243] = 106;
        test_data[2243] = 33'd8183296017;
        test_addr[2244] = 437;
        test_data[2244] = 33'd6784118135;
        test_addr[2245] = 254;
        test_data[2245] = 33'd8533089254;
        test_addr[2246] = 751;
        test_data[2246] = 33'd2723074538;
        test_addr[2247] = 969;
        test_data[2247] = 33'd1632363957;
        test_addr[2248] = 167;
        test_data[2248] = 33'd188544578;
        test_addr[2249] = 511;
        test_data[2249] = 33'd308446067;
        test_addr[2250] = 56;
        test_data[2250] = 33'd3847507083;
        test_addr[2251] = 828;
        test_data[2251] = 33'd2346462542;
        test_addr[2252] = 372;
        test_data[2252] = 33'd3706783982;
        test_addr[2253] = 8;
        test_data[2253] = 33'd5773335490;
        test_addr[2254] = 1020;
        test_data[2254] = 33'd1993492834;
        test_addr[2255] = 676;
        test_data[2255] = 33'd1174454579;
        test_addr[2256] = 145;
        test_data[2256] = 33'd5509182353;
        test_addr[2257] = 536;
        test_data[2257] = 33'd1677816877;
        test_addr[2258] = 384;
        test_data[2258] = 33'd7070588422;
        test_addr[2259] = 213;
        test_data[2259] = 33'd2155161093;
        test_addr[2260] = 503;
        test_data[2260] = 33'd7922472969;
        test_addr[2261] = 348;
        test_data[2261] = 33'd3222427471;
        test_addr[2262] = 390;
        test_data[2262] = 33'd909123417;
        test_addr[2263] = 541;
        test_data[2263] = 33'd4208840303;
        test_addr[2264] = 85;
        test_data[2264] = 33'd3303270017;
        test_addr[2265] = 846;
        test_data[2265] = 33'd4626776678;
        test_addr[2266] = 136;
        test_data[2266] = 33'd8215380217;
        test_addr[2267] = 1004;
        test_data[2267] = 33'd8136772519;
        test_addr[2268] = 658;
        test_data[2268] = 33'd8582733612;
        test_addr[2269] = 328;
        test_data[2269] = 33'd5319566575;
        test_addr[2270] = 885;
        test_data[2270] = 33'd728215166;
        test_addr[2271] = 334;
        test_data[2271] = 33'd3431054307;
        test_addr[2272] = 853;
        test_data[2272] = 33'd3599534504;
        test_addr[2273] = 727;
        test_data[2273] = 33'd4061007751;
        test_addr[2274] = 935;
        test_data[2274] = 33'd3858261570;
        test_addr[2275] = 658;
        test_data[2275] = 33'd4930166811;
        test_addr[2276] = 437;
        test_data[2276] = 33'd2489150839;
        test_addr[2277] = 18;
        test_data[2277] = 33'd3370794791;
        test_addr[2278] = 866;
        test_data[2278] = 33'd6881866486;
        test_addr[2279] = 897;
        test_data[2279] = 33'd4543160669;
        test_addr[2280] = 615;
        test_data[2280] = 33'd2136755942;
        test_addr[2281] = 926;
        test_data[2281] = 33'd7817684517;
        test_addr[2282] = 41;
        test_data[2282] = 33'd1738554561;
        test_addr[2283] = 788;
        test_data[2283] = 33'd3121816568;
        test_addr[2284] = 82;
        test_data[2284] = 33'd1180769850;
        test_addr[2285] = 818;
        test_data[2285] = 33'd702408417;
        test_addr[2286] = 467;
        test_data[2286] = 33'd5537426286;
        test_addr[2287] = 219;
        test_data[2287] = 33'd308900539;
        test_addr[2288] = 712;
        test_data[2288] = 33'd7601294151;
        test_addr[2289] = 889;
        test_data[2289] = 33'd4420085022;
        test_addr[2290] = 766;
        test_data[2290] = 33'd1804301512;
        test_addr[2291] = 790;
        test_data[2291] = 33'd3048710191;
        test_addr[2292] = 989;
        test_data[2292] = 33'd4492828763;
        test_addr[2293] = 875;
        test_data[2293] = 33'd5037940627;
        test_addr[2294] = 601;
        test_data[2294] = 33'd2919076942;
        test_addr[2295] = 738;
        test_data[2295] = 33'd5136843289;
        test_addr[2296] = 649;
        test_data[2296] = 33'd6427719060;
        test_addr[2297] = 697;
        test_data[2297] = 33'd3089205481;
        test_addr[2298] = 904;
        test_data[2298] = 33'd580095324;
        test_addr[2299] = 584;
        test_data[2299] = 33'd5354288876;
        test_addr[2300] = 116;
        test_data[2300] = 33'd920627105;
        test_addr[2301] = 295;
        test_data[2301] = 33'd7489464297;
        test_addr[2302] = 230;
        test_data[2302] = 33'd3123327297;
        test_addr[2303] = 880;
        test_data[2303] = 33'd2124676183;
        test_addr[2304] = 953;
        test_data[2304] = 33'd1370236496;
        test_addr[2305] = 770;
        test_data[2305] = 33'd3253604653;
        test_addr[2306] = 452;
        test_data[2306] = 33'd4495689235;
        test_addr[2307] = 89;
        test_data[2307] = 33'd4495969493;
        test_addr[2308] = 955;
        test_data[2308] = 33'd199830729;
        test_addr[2309] = 249;
        test_data[2309] = 33'd3994305534;
        test_addr[2310] = 875;
        test_data[2310] = 33'd6587307734;
        test_addr[2311] = 637;
        test_data[2311] = 33'd1672692856;
        test_addr[2312] = 291;
        test_data[2312] = 33'd4323708592;
        test_addr[2313] = 318;
        test_data[2313] = 33'd1218864492;
        test_addr[2314] = 624;
        test_data[2314] = 33'd5159297085;
        test_addr[2315] = 169;
        test_data[2315] = 33'd1816155489;
        test_addr[2316] = 34;
        test_data[2316] = 33'd7471832863;
        test_addr[2317] = 923;
        test_data[2317] = 33'd2479546912;
        test_addr[2318] = 272;
        test_data[2318] = 33'd478200901;
        test_addr[2319] = 821;
        test_data[2319] = 33'd1331449937;
        test_addr[2320] = 365;
        test_data[2320] = 33'd369210451;
        test_addr[2321] = 709;
        test_data[2321] = 33'd1267071129;
        test_addr[2322] = 275;
        test_data[2322] = 33'd4044162456;
        test_addr[2323] = 322;
        test_data[2323] = 33'd3243207308;
        test_addr[2324] = 902;
        test_data[2324] = 33'd6667354578;
        test_addr[2325] = 764;
        test_data[2325] = 33'd82671605;
        test_addr[2326] = 683;
        test_data[2326] = 33'd6328370987;
        test_addr[2327] = 318;
        test_data[2327] = 33'd1218864492;
        test_addr[2328] = 776;
        test_data[2328] = 33'd769284591;
        test_addr[2329] = 706;
        test_data[2329] = 33'd785242298;
        test_addr[2330] = 522;
        test_data[2330] = 33'd4304962878;
        test_addr[2331] = 342;
        test_data[2331] = 33'd1814882452;
        test_addr[2332] = 390;
        test_data[2332] = 33'd909123417;
        test_addr[2333] = 1006;
        test_data[2333] = 33'd2390501042;
        test_addr[2334] = 872;
        test_data[2334] = 33'd3871519302;
        test_addr[2335] = 900;
        test_data[2335] = 33'd3715729542;
        test_addr[2336] = 64;
        test_data[2336] = 33'd3038722049;
        test_addr[2337] = 275;
        test_data[2337] = 33'd8165126272;
        test_addr[2338] = 857;
        test_data[2338] = 33'd1320604479;
        test_addr[2339] = 680;
        test_data[2339] = 33'd8402810508;
        test_addr[2340] = 130;
        test_data[2340] = 33'd1268433295;
        test_addr[2341] = 431;
        test_data[2341] = 33'd7722785918;
        test_addr[2342] = 261;
        test_data[2342] = 33'd4668518653;
        test_addr[2343] = 847;
        test_data[2343] = 33'd196428976;
        test_addr[2344] = 566;
        test_data[2344] = 33'd3593853367;
        test_addr[2345] = 465;
        test_data[2345] = 33'd896820312;
        test_addr[2346] = 228;
        test_data[2346] = 33'd4827997493;
        test_addr[2347] = 1;
        test_data[2347] = 33'd2545176946;
        test_addr[2348] = 234;
        test_data[2348] = 33'd3874139594;
        test_addr[2349] = 886;
        test_data[2349] = 33'd7256702761;
        test_addr[2350] = 611;
        test_data[2350] = 33'd803685859;
        test_addr[2351] = 427;
        test_data[2351] = 33'd3998550133;
        test_addr[2352] = 890;
        test_data[2352] = 33'd2018427355;
        test_addr[2353] = 488;
        test_data[2353] = 33'd839680804;
        test_addr[2354] = 385;
        test_data[2354] = 33'd7242686252;
        test_addr[2355] = 565;
        test_data[2355] = 33'd7890552546;
        test_addr[2356] = 265;
        test_data[2356] = 33'd3802763157;
        test_addr[2357] = 755;
        test_data[2357] = 33'd2070820228;
        test_addr[2358] = 1010;
        test_data[2358] = 33'd4501859999;
        test_addr[2359] = 223;
        test_data[2359] = 33'd3210078290;
        test_addr[2360] = 1001;
        test_data[2360] = 33'd7308170596;
        test_addr[2361] = 542;
        test_data[2361] = 33'd2688370830;
        test_addr[2362] = 344;
        test_data[2362] = 33'd6694505707;
        test_addr[2363] = 611;
        test_data[2363] = 33'd8235616715;
        test_addr[2364] = 879;
        test_data[2364] = 33'd2227416794;
        test_addr[2365] = 563;
        test_data[2365] = 33'd4151707470;
        test_addr[2366] = 144;
        test_data[2366] = 33'd4214779887;
        test_addr[2367] = 103;
        test_data[2367] = 33'd7808076481;
        test_addr[2368] = 973;
        test_data[2368] = 33'd986805218;
        test_addr[2369] = 836;
        test_data[2369] = 33'd1052769268;
        test_addr[2370] = 972;
        test_data[2370] = 33'd7045577130;
        test_addr[2371] = 196;
        test_data[2371] = 33'd6086400782;
        test_addr[2372] = 364;
        test_data[2372] = 33'd4222053268;
        test_addr[2373] = 360;
        test_data[2373] = 33'd40490138;
        test_addr[2374] = 437;
        test_data[2374] = 33'd2489150839;
        test_addr[2375] = 855;
        test_data[2375] = 33'd4608367523;
        test_addr[2376] = 661;
        test_data[2376] = 33'd7562028680;
        test_addr[2377] = 155;
        test_data[2377] = 33'd6920961997;
        test_addr[2378] = 982;
        test_data[2378] = 33'd3029117888;
        test_addr[2379] = 859;
        test_data[2379] = 33'd1314706587;
        test_addr[2380] = 801;
        test_data[2380] = 33'd448058807;
        test_addr[2381] = 68;
        test_data[2381] = 33'd2031775880;
        test_addr[2382] = 479;
        test_data[2382] = 33'd3763673002;
        test_addr[2383] = 61;
        test_data[2383] = 33'd8506161349;
        test_addr[2384] = 179;
        test_data[2384] = 33'd3433493149;
        test_addr[2385] = 976;
        test_data[2385] = 33'd3839524366;
        test_addr[2386] = 448;
        test_data[2386] = 33'd2388061351;
        test_addr[2387] = 897;
        test_data[2387] = 33'd4909155405;
        test_addr[2388] = 153;
        test_data[2388] = 33'd632865373;
        test_addr[2389] = 942;
        test_data[2389] = 33'd2133741656;
        test_addr[2390] = 130;
        test_data[2390] = 33'd5117731653;
        test_addr[2391] = 843;
        test_data[2391] = 33'd5560499837;
        test_addr[2392] = 834;
        test_data[2392] = 33'd7720126015;
        test_addr[2393] = 733;
        test_data[2393] = 33'd8214366487;
        test_addr[2394] = 313;
        test_data[2394] = 33'd2105637580;
        test_addr[2395] = 113;
        test_data[2395] = 33'd2029943915;
        test_addr[2396] = 113;
        test_data[2396] = 33'd2029943915;
        test_addr[2397] = 262;
        test_data[2397] = 33'd3966004824;
        test_addr[2398] = 244;
        test_data[2398] = 33'd656960195;
        test_addr[2399] = 1006;
        test_data[2399] = 33'd2390501042;
        test_addr[2400] = 591;
        test_data[2400] = 33'd3406733999;
        test_addr[2401] = 435;
        test_data[2401] = 33'd3843532341;
        test_addr[2402] = 735;
        test_data[2402] = 33'd1228527252;
        test_addr[2403] = 628;
        test_data[2403] = 33'd3902713659;
        test_addr[2404] = 796;
        test_data[2404] = 33'd6145444028;
        test_addr[2405] = 580;
        test_data[2405] = 33'd4568718784;
        test_addr[2406] = 596;
        test_data[2406] = 33'd4087896024;
        test_addr[2407] = 92;
        test_data[2407] = 33'd5180956050;
        test_addr[2408] = 180;
        test_data[2408] = 33'd4026446541;
        test_addr[2409] = 238;
        test_data[2409] = 33'd291352294;
        test_addr[2410] = 737;
        test_data[2410] = 33'd4499394865;
        test_addr[2411] = 612;
        test_data[2411] = 33'd4539353342;
        test_addr[2412] = 23;
        test_data[2412] = 33'd1087399442;
        test_addr[2413] = 386;
        test_data[2413] = 33'd5426199134;
        test_addr[2414] = 131;
        test_data[2414] = 33'd813280569;
        test_addr[2415] = 137;
        test_data[2415] = 33'd3806722747;
        test_addr[2416] = 404;
        test_data[2416] = 33'd7526840985;
        test_addr[2417] = 683;
        test_data[2417] = 33'd2033403691;
        test_addr[2418] = 973;
        test_data[2418] = 33'd986805218;
        test_addr[2419] = 847;
        test_data[2419] = 33'd196428976;
        test_addr[2420] = 282;
        test_data[2420] = 33'd5502154964;
        test_addr[2421] = 778;
        test_data[2421] = 33'd6623421118;
        test_addr[2422] = 885;
        test_data[2422] = 33'd7992909893;
        test_addr[2423] = 959;
        test_data[2423] = 33'd910132403;
        test_addr[2424] = 103;
        test_data[2424] = 33'd7218880973;
        test_addr[2425] = 413;
        test_data[2425] = 33'd3563808226;
        test_addr[2426] = 704;
        test_data[2426] = 33'd7891837135;
        test_addr[2427] = 428;
        test_data[2427] = 33'd1801007473;
        test_addr[2428] = 560;
        test_data[2428] = 33'd3890402307;
        test_addr[2429] = 271;
        test_data[2429] = 33'd644631020;
        test_addr[2430] = 0;
        test_data[2430] = 33'd5881492295;
        test_addr[2431] = 404;
        test_data[2431] = 33'd3231873689;
        test_addr[2432] = 707;
        test_data[2432] = 33'd6389108407;
        test_addr[2433] = 136;
        test_data[2433] = 33'd3920412921;
        test_addr[2434] = 266;
        test_data[2434] = 33'd398595192;
        test_addr[2435] = 16;
        test_data[2435] = 33'd2233696814;
        test_addr[2436] = 612;
        test_data[2436] = 33'd244386046;
        test_addr[2437] = 45;
        test_data[2437] = 33'd5074297821;
        test_addr[2438] = 784;
        test_data[2438] = 33'd5060732098;
        test_addr[2439] = 602;
        test_data[2439] = 33'd3481104526;
        test_addr[2440] = 198;
        test_data[2440] = 33'd1601624005;
        test_addr[2441] = 362;
        test_data[2441] = 33'd4225808861;
        test_addr[2442] = 255;
        test_data[2442] = 33'd1916824779;
        test_addr[2443] = 692;
        test_data[2443] = 33'd6148442540;
        test_addr[2444] = 717;
        test_data[2444] = 33'd3881300217;
        test_addr[2445] = 933;
        test_data[2445] = 33'd2246106299;
        test_addr[2446] = 97;
        test_data[2446] = 33'd1378927735;
        test_addr[2447] = 985;
        test_data[2447] = 33'd2974518957;
        test_addr[2448] = 652;
        test_data[2448] = 33'd7810425231;
        test_addr[2449] = 100;
        test_data[2449] = 33'd4815712175;
        test_addr[2450] = 274;
        test_data[2450] = 33'd190441195;
        test_addr[2451] = 948;
        test_data[2451] = 33'd1756278281;
        test_addr[2452] = 52;
        test_data[2452] = 33'd3594104512;
        test_addr[2453] = 789;
        test_data[2453] = 33'd2899379877;
        test_addr[2454] = 630;
        test_data[2454] = 33'd142622312;
        test_addr[2455] = 734;
        test_data[2455] = 33'd3464739256;
        test_addr[2456] = 470;
        test_data[2456] = 33'd408988608;
        test_addr[2457] = 673;
        test_data[2457] = 33'd41814705;
        test_addr[2458] = 98;
        test_data[2458] = 33'd6500919089;
        test_addr[2459] = 426;
        test_data[2459] = 33'd7208989612;
        test_addr[2460] = 709;
        test_data[2460] = 33'd7656830057;
        test_addr[2461] = 455;
        test_data[2461] = 33'd2867352729;
        test_addr[2462] = 44;
        test_data[2462] = 33'd8565640083;
        test_addr[2463] = 598;
        test_data[2463] = 33'd3684002157;
        test_addr[2464] = 777;
        test_data[2464] = 33'd1706937674;
        test_addr[2465] = 889;
        test_data[2465] = 33'd125117726;
        test_addr[2466] = 409;
        test_data[2466] = 33'd1313692123;
        test_addr[2467] = 579;
        test_data[2467] = 33'd2718604588;
        test_addr[2468] = 58;
        test_data[2468] = 33'd463636514;
        test_addr[2469] = 295;
        test_data[2469] = 33'd5008262652;
        test_addr[2470] = 797;
        test_data[2470] = 33'd8086720465;
        test_addr[2471] = 354;
        test_data[2471] = 33'd6601391683;
        test_addr[2472] = 872;
        test_data[2472] = 33'd8329920513;
        test_addr[2473] = 861;
        test_data[2473] = 33'd3320468775;
        test_addr[2474] = 217;
        test_data[2474] = 33'd3904384728;
        test_addr[2475] = 436;
        test_data[2475] = 33'd7058285698;
        test_addr[2476] = 540;
        test_data[2476] = 33'd8252533019;
        test_addr[2477] = 911;
        test_data[2477] = 33'd2047098942;
        test_addr[2478] = 460;
        test_data[2478] = 33'd1546315615;
        test_addr[2479] = 994;
        test_data[2479] = 33'd4477219491;
        test_addr[2480] = 838;
        test_data[2480] = 33'd1113939390;
        test_addr[2481] = 445;
        test_data[2481] = 33'd550922961;
        test_addr[2482] = 549;
        test_data[2482] = 33'd5599632497;
        test_addr[2483] = 200;
        test_data[2483] = 33'd4007449550;
        test_addr[2484] = 302;
        test_data[2484] = 33'd6505288025;
        test_addr[2485] = 150;
        test_data[2485] = 33'd735908553;
        test_addr[2486] = 72;
        test_data[2486] = 33'd7127641884;
        test_addr[2487] = 717;
        test_data[2487] = 33'd4404868719;
        test_addr[2488] = 363;
        test_data[2488] = 33'd2998056081;
        test_addr[2489] = 788;
        test_data[2489] = 33'd3121816568;
        test_addr[2490] = 113;
        test_data[2490] = 33'd2029943915;
        test_addr[2491] = 142;
        test_data[2491] = 33'd2983160463;
        test_addr[2492] = 446;
        test_data[2492] = 33'd1909467616;
        test_addr[2493] = 730;
        test_data[2493] = 33'd363081077;
        test_addr[2494] = 658;
        test_data[2494] = 33'd635199515;
        test_addr[2495] = 64;
        test_data[2495] = 33'd3038722049;
        test_addr[2496] = 835;
        test_data[2496] = 33'd2129932696;
        test_addr[2497] = 662;
        test_data[2497] = 33'd4677729244;
        test_addr[2498] = 107;
        test_data[2498] = 33'd4243198286;
        test_addr[2499] = 975;
        test_data[2499] = 33'd1686953869;
        test_addr[2500] = 821;
        test_data[2500] = 33'd5968904785;
        test_addr[2501] = 714;
        test_data[2501] = 33'd761390289;
        test_addr[2502] = 102;
        test_data[2502] = 33'd1124317209;
        test_addr[2503] = 76;
        test_data[2503] = 33'd8074482355;
        test_addr[2504] = 986;
        test_data[2504] = 33'd2081595685;
        test_addr[2505] = 836;
        test_data[2505] = 33'd1052769268;
        test_addr[2506] = 580;
        test_data[2506] = 33'd6602941603;
        test_addr[2507] = 782;
        test_data[2507] = 33'd4948194028;
        test_addr[2508] = 600;
        test_data[2508] = 33'd1402039586;
        test_addr[2509] = 310;
        test_data[2509] = 33'd3692301779;
        test_addr[2510] = 144;
        test_data[2510] = 33'd4214779887;
        test_addr[2511] = 876;
        test_data[2511] = 33'd7077828655;
        test_addr[2512] = 356;
        test_data[2512] = 33'd6600338461;
        test_addr[2513] = 724;
        test_data[2513] = 33'd4230629022;
        test_addr[2514] = 1012;
        test_data[2514] = 33'd4031553092;
        test_addr[2515] = 890;
        test_data[2515] = 33'd6791844085;
        test_addr[2516] = 697;
        test_data[2516] = 33'd5438101706;
        test_addr[2517] = 87;
        test_data[2517] = 33'd6977262976;
        test_addr[2518] = 688;
        test_data[2518] = 33'd7143529981;
        test_addr[2519] = 714;
        test_data[2519] = 33'd761390289;
        test_addr[2520] = 245;
        test_data[2520] = 33'd7624746068;
        test_addr[2521] = 35;
        test_data[2521] = 33'd6620224688;
        test_addr[2522] = 327;
        test_data[2522] = 33'd2012735954;
        test_addr[2523] = 962;
        test_data[2523] = 33'd6588613504;
        test_addr[2524] = 311;
        test_data[2524] = 33'd3503918147;
        test_addr[2525] = 246;
        test_data[2525] = 33'd1635138116;
        test_addr[2526] = 556;
        test_data[2526] = 33'd4599692122;
        test_addr[2527] = 696;
        test_data[2527] = 33'd2694337344;
        test_addr[2528] = 694;
        test_data[2528] = 33'd4915529711;
        test_addr[2529] = 954;
        test_data[2529] = 33'd1594670622;
        test_addr[2530] = 328;
        test_data[2530] = 33'd1024599279;
        test_addr[2531] = 699;
        test_data[2531] = 33'd5435045928;
        test_addr[2532] = 786;
        test_data[2532] = 33'd2790845645;
        test_addr[2533] = 266;
        test_data[2533] = 33'd7279864570;
        test_addr[2534] = 397;
        test_data[2534] = 33'd5007129743;
        test_addr[2535] = 475;
        test_data[2535] = 33'd6703834173;
        test_addr[2536] = 109;
        test_data[2536] = 33'd6921059266;
        test_addr[2537] = 951;
        test_data[2537] = 33'd511634929;
        test_addr[2538] = 18;
        test_data[2538] = 33'd3370794791;
        test_addr[2539] = 492;
        test_data[2539] = 33'd7175142947;
        test_addr[2540] = 722;
        test_data[2540] = 33'd8160917662;
        test_addr[2541] = 775;
        test_data[2541] = 33'd4264175710;
        test_addr[2542] = 337;
        test_data[2542] = 33'd7087052729;
        test_addr[2543] = 686;
        test_data[2543] = 33'd318457616;
        test_addr[2544] = 282;
        test_data[2544] = 33'd5568603449;
        test_addr[2545] = 666;
        test_data[2545] = 33'd4838698039;
        test_addr[2546] = 983;
        test_data[2546] = 33'd509354105;
        test_addr[2547] = 450;
        test_data[2547] = 33'd2461350224;
        test_addr[2548] = 617;
        test_data[2548] = 33'd883935601;
        test_addr[2549] = 82;
        test_data[2549] = 33'd1180769850;
        test_addr[2550] = 789;
        test_data[2550] = 33'd2899379877;
        test_addr[2551] = 374;
        test_data[2551] = 33'd2011634502;
        test_addr[2552] = 121;
        test_data[2552] = 33'd157354656;
        test_addr[2553] = 381;
        test_data[2553] = 33'd1838811245;
        test_addr[2554] = 111;
        test_data[2554] = 33'd3462749259;
        test_addr[2555] = 664;
        test_data[2555] = 33'd1694872111;
        test_addr[2556] = 433;
        test_data[2556] = 33'd5561069201;
        test_addr[2557] = 343;
        test_data[2557] = 33'd6744936583;
        test_addr[2558] = 274;
        test_data[2558] = 33'd190441195;
        test_addr[2559] = 250;
        test_data[2559] = 33'd6228569223;
        test_addr[2560] = 3;
        test_data[2560] = 33'd24445434;
        test_addr[2561] = 406;
        test_data[2561] = 33'd1667658830;
        test_addr[2562] = 434;
        test_data[2562] = 33'd188263586;
        test_addr[2563] = 104;
        test_data[2563] = 33'd6303654149;
        test_addr[2564] = 950;
        test_data[2564] = 33'd478080935;
        test_addr[2565] = 645;
        test_data[2565] = 33'd543326322;
        test_addr[2566] = 541;
        test_data[2566] = 33'd4208840303;
        test_addr[2567] = 470;
        test_data[2567] = 33'd408988608;
        test_addr[2568] = 394;
        test_data[2568] = 33'd6151588535;
        test_addr[2569] = 868;
        test_data[2569] = 33'd5887100844;
        test_addr[2570] = 955;
        test_data[2570] = 33'd6621034010;
        test_addr[2571] = 651;
        test_data[2571] = 33'd2210885566;
        test_addr[2572] = 845;
        test_data[2572] = 33'd1963746399;
        test_addr[2573] = 362;
        test_data[2573] = 33'd8033338721;
        test_addr[2574] = 848;
        test_data[2574] = 33'd5403081423;
        test_addr[2575] = 736;
        test_data[2575] = 33'd1931613996;
        test_addr[2576] = 895;
        test_data[2576] = 33'd7465816292;
        test_addr[2577] = 453;
        test_data[2577] = 33'd2561706829;
        test_addr[2578] = 205;
        test_data[2578] = 33'd6215367386;
        test_addr[2579] = 135;
        test_data[2579] = 33'd69857205;
        test_addr[2580] = 712;
        test_data[2580] = 33'd6550650315;
        test_addr[2581] = 737;
        test_data[2581] = 33'd5946931738;
        test_addr[2582] = 716;
        test_data[2582] = 33'd3103417907;
        test_addr[2583] = 401;
        test_data[2583] = 33'd2799343604;
        test_addr[2584] = 553;
        test_data[2584] = 33'd7019763371;
        test_addr[2585] = 902;
        test_data[2585] = 33'd2372387282;
        test_addr[2586] = 8;
        test_data[2586] = 33'd1478368194;
        test_addr[2587] = 830;
        test_data[2587] = 33'd6903434084;
        test_addr[2588] = 219;
        test_data[2588] = 33'd8471635372;
        test_addr[2589] = 538;
        test_data[2589] = 33'd4321225144;
        test_addr[2590] = 503;
        test_data[2590] = 33'd5486440831;
        test_addr[2591] = 273;
        test_data[2591] = 33'd56693191;
        test_addr[2592] = 197;
        test_data[2592] = 33'd2393364357;
        test_addr[2593] = 61;
        test_data[2593] = 33'd4211194053;
        test_addr[2594] = 869;
        test_data[2594] = 33'd2336492666;
        test_addr[2595] = 768;
        test_data[2595] = 33'd8006448719;
        test_addr[2596] = 416;
        test_data[2596] = 33'd3819993292;
        test_addr[2597] = 880;
        test_data[2597] = 33'd2124676183;
        test_addr[2598] = 328;
        test_data[2598] = 33'd6004527447;
        test_addr[2599] = 292;
        test_data[2599] = 33'd2819396262;
        test_addr[2600] = 643;
        test_data[2600] = 33'd6129206424;
        test_addr[2601] = 990;
        test_data[2601] = 33'd4082014275;
        test_addr[2602] = 942;
        test_data[2602] = 33'd2133741656;
        test_addr[2603] = 665;
        test_data[2603] = 33'd1128756264;
        test_addr[2604] = 457;
        test_data[2604] = 33'd6320375093;
        test_addr[2605] = 135;
        test_data[2605] = 33'd69857205;
        test_addr[2606] = 930;
        test_data[2606] = 33'd2007557742;
        test_addr[2607] = 757;
        test_data[2607] = 33'd7023070098;
        test_addr[2608] = 489;
        test_data[2608] = 33'd3603165913;
        test_addr[2609] = 81;
        test_data[2609] = 33'd3391775223;
        test_addr[2610] = 629;
        test_data[2610] = 33'd1773980868;
        test_addr[2611] = 903;
        test_data[2611] = 33'd4854858965;
        test_addr[2612] = 596;
        test_data[2612] = 33'd5967439355;
        test_addr[2613] = 156;
        test_data[2613] = 33'd3852022963;
        test_addr[2614] = 159;
        test_data[2614] = 33'd571794251;
        test_addr[2615] = 95;
        test_data[2615] = 33'd7522062609;
        test_addr[2616] = 529;
        test_data[2616] = 33'd4702799624;
        test_addr[2617] = 416;
        test_data[2617] = 33'd3819993292;
        test_addr[2618] = 33;
        test_data[2618] = 33'd1484688907;
        test_addr[2619] = 261;
        test_data[2619] = 33'd7160722995;
        test_addr[2620] = 946;
        test_data[2620] = 33'd1789457252;
        test_addr[2621] = 290;
        test_data[2621] = 33'd3989670362;
        test_addr[2622] = 74;
        test_data[2622] = 33'd3405503829;
        test_addr[2623] = 661;
        test_data[2623] = 33'd3267061384;
        test_addr[2624] = 425;
        test_data[2624] = 33'd6527801575;
        test_addr[2625] = 27;
        test_data[2625] = 33'd4678896834;
        test_addr[2626] = 448;
        test_data[2626] = 33'd2388061351;
        test_addr[2627] = 438;
        test_data[2627] = 33'd2860390341;
        test_addr[2628] = 124;
        test_data[2628] = 33'd7637667207;
        test_addr[2629] = 264;
        test_data[2629] = 33'd687477629;
        test_addr[2630] = 916;
        test_data[2630] = 33'd1736915697;
        test_addr[2631] = 660;
        test_data[2631] = 33'd1826723096;
        test_addr[2632] = 796;
        test_data[2632] = 33'd6743054685;
        test_addr[2633] = 285;
        test_data[2633] = 33'd1566790510;
        test_addr[2634] = 814;
        test_data[2634] = 33'd662516995;
        test_addr[2635] = 826;
        test_data[2635] = 33'd690145171;
        test_addr[2636] = 884;
        test_data[2636] = 33'd5794233438;
        test_addr[2637] = 229;
        test_data[2637] = 33'd920626449;
        test_addr[2638] = 456;
        test_data[2638] = 33'd7330508917;
        test_addr[2639] = 580;
        test_data[2639] = 33'd2307974307;
        test_addr[2640] = 557;
        test_data[2640] = 33'd4627833013;
        test_addr[2641] = 1004;
        test_data[2641] = 33'd6068961283;
        test_addr[2642] = 922;
        test_data[2642] = 33'd715587172;
        test_addr[2643] = 49;
        test_data[2643] = 33'd751512591;
        test_addr[2644] = 743;
        test_data[2644] = 33'd3612336317;
        test_addr[2645] = 335;
        test_data[2645] = 33'd2081762056;
        test_addr[2646] = 143;
        test_data[2646] = 33'd796190208;
        test_addr[2647] = 757;
        test_data[2647] = 33'd4502169927;
        test_addr[2648] = 222;
        test_data[2648] = 33'd3784662317;
        test_addr[2649] = 838;
        test_data[2649] = 33'd1113939390;
        test_addr[2650] = 97;
        test_data[2650] = 33'd1378927735;
        test_addr[2651] = 907;
        test_data[2651] = 33'd4168846095;
        test_addr[2652] = 725;
        test_data[2652] = 33'd1347397057;
        test_addr[2653] = 6;
        test_data[2653] = 33'd1280683540;
        test_addr[2654] = 317;
        test_data[2654] = 33'd6879706816;
        test_addr[2655] = 157;
        test_data[2655] = 33'd5929256640;
        test_addr[2656] = 780;
        test_data[2656] = 33'd404411201;
        test_addr[2657] = 418;
        test_data[2657] = 33'd6723766007;
        test_addr[2658] = 591;
        test_data[2658] = 33'd7021289310;
        test_addr[2659] = 599;
        test_data[2659] = 33'd4446249921;
        test_addr[2660] = 856;
        test_data[2660] = 33'd975862316;
        test_addr[2661] = 607;
        test_data[2661] = 33'd6147980072;
        test_addr[2662] = 735;
        test_data[2662] = 33'd4699784797;
        test_addr[2663] = 823;
        test_data[2663] = 33'd1932951958;
        test_addr[2664] = 613;
        test_data[2664] = 33'd8559343628;
        test_addr[2665] = 518;
        test_data[2665] = 33'd2506176115;
        test_addr[2666] = 749;
        test_data[2666] = 33'd987435852;
        test_addr[2667] = 247;
        test_data[2667] = 33'd4009011063;
        test_addr[2668] = 883;
        test_data[2668] = 33'd1795705404;
        test_addr[2669] = 633;
        test_data[2669] = 33'd7255536440;
        test_addr[2670] = 366;
        test_data[2670] = 33'd7167074511;
        test_addr[2671] = 315;
        test_data[2671] = 33'd3577492034;
        test_addr[2672] = 558;
        test_data[2672] = 33'd8482512041;
        test_addr[2673] = 931;
        test_data[2673] = 33'd2803979244;
        test_addr[2674] = 402;
        test_data[2674] = 33'd1208032225;
        test_addr[2675] = 506;
        test_data[2675] = 33'd3145293850;
        test_addr[2676] = 997;
        test_data[2676] = 33'd7522627152;
        test_addr[2677] = 674;
        test_data[2677] = 33'd6438688497;
        test_addr[2678] = 221;
        test_data[2678] = 33'd720358563;
        test_addr[2679] = 365;
        test_data[2679] = 33'd369210451;
        test_addr[2680] = 543;
        test_data[2680] = 33'd3369326361;
        test_addr[2681] = 300;
        test_data[2681] = 33'd532524759;
        test_addr[2682] = 668;
        test_data[2682] = 33'd6589462861;
        test_addr[2683] = 18;
        test_data[2683] = 33'd3370794791;
        test_addr[2684] = 659;
        test_data[2684] = 33'd7882082485;
        test_addr[2685] = 428;
        test_data[2685] = 33'd1801007473;
        test_addr[2686] = 659;
        test_data[2686] = 33'd8588020703;
        test_addr[2687] = 528;
        test_data[2687] = 33'd3661790944;
        test_addr[2688] = 818;
        test_data[2688] = 33'd6354211875;
        test_addr[2689] = 169;
        test_data[2689] = 33'd6171954597;
        test_addr[2690] = 504;
        test_data[2690] = 33'd2373341895;
        test_addr[2691] = 419;
        test_data[2691] = 33'd4133168253;
        test_addr[2692] = 644;
        test_data[2692] = 33'd3810663823;
        test_addr[2693] = 562;
        test_data[2693] = 33'd579089702;
        test_addr[2694] = 820;
        test_data[2694] = 33'd4175331955;
        test_addr[2695] = 163;
        test_data[2695] = 33'd2222230867;
        test_addr[2696] = 961;
        test_data[2696] = 33'd2071565022;
        test_addr[2697] = 103;
        test_data[2697] = 33'd2923913677;
        test_addr[2698] = 144;
        test_data[2698] = 33'd4214779887;
        test_addr[2699] = 776;
        test_data[2699] = 33'd769284591;
        test_addr[2700] = 18;
        test_data[2700] = 33'd6312308070;
        test_addr[2701] = 273;
        test_data[2701] = 33'd56693191;
        test_addr[2702] = 724;
        test_data[2702] = 33'd4230629022;
        test_addr[2703] = 736;
        test_data[2703] = 33'd6899190917;
        test_addr[2704] = 607;
        test_data[2704] = 33'd1853012776;
        test_addr[2705] = 367;
        test_data[2705] = 33'd1561819636;
        test_addr[2706] = 228;
        test_data[2706] = 33'd533030197;
        test_addr[2707] = 993;
        test_data[2707] = 33'd2909818976;
        test_addr[2708] = 880;
        test_data[2708] = 33'd2124676183;
        test_addr[2709] = 147;
        test_data[2709] = 33'd2764225137;
        test_addr[2710] = 47;
        test_data[2710] = 33'd1684233673;
        test_addr[2711] = 516;
        test_data[2711] = 33'd3235422805;
        test_addr[2712] = 187;
        test_data[2712] = 33'd3002320632;
        test_addr[2713] = 846;
        test_data[2713] = 33'd331809382;
        test_addr[2714] = 777;
        test_data[2714] = 33'd7551810475;
        test_addr[2715] = 306;
        test_data[2715] = 33'd1818292495;
        test_addr[2716] = 879;
        test_data[2716] = 33'd2227416794;
        test_addr[2717] = 984;
        test_data[2717] = 33'd3168600535;
        test_addr[2718] = 804;
        test_data[2718] = 33'd2469310094;
        test_addr[2719] = 247;
        test_data[2719] = 33'd4009011063;
        test_addr[2720] = 1023;
        test_data[2720] = 33'd7681764131;
        test_addr[2721] = 622;
        test_data[2721] = 33'd5546579813;
        test_addr[2722] = 462;
        test_data[2722] = 33'd6947911624;
        test_addr[2723] = 908;
        test_data[2723] = 33'd1704854364;
        test_addr[2724] = 777;
        test_data[2724] = 33'd3256843179;
        test_addr[2725] = 952;
        test_data[2725] = 33'd4073189063;
        test_addr[2726] = 388;
        test_data[2726] = 33'd800990285;
        test_addr[2727] = 890;
        test_data[2727] = 33'd2496876789;
        test_addr[2728] = 812;
        test_data[2728] = 33'd1111087967;
        test_addr[2729] = 403;
        test_data[2729] = 33'd2351946442;
        test_addr[2730] = 192;
        test_data[2730] = 33'd2694434016;
        test_addr[2731] = 196;
        test_data[2731] = 33'd1791433486;
        test_addr[2732] = 932;
        test_data[2732] = 33'd4275128377;
        test_addr[2733] = 110;
        test_data[2733] = 33'd6258519054;
        test_addr[2734] = 174;
        test_data[2734] = 33'd3604100316;
        test_addr[2735] = 137;
        test_data[2735] = 33'd3806722747;
        test_addr[2736] = 151;
        test_data[2736] = 33'd2126478811;
        test_addr[2737] = 247;
        test_data[2737] = 33'd4009011063;
        test_addr[2738] = 632;
        test_data[2738] = 33'd162213990;
        test_addr[2739] = 119;
        test_data[2739] = 33'd2763234325;
        test_addr[2740] = 823;
        test_data[2740] = 33'd1932951958;
        test_addr[2741] = 872;
        test_data[2741] = 33'd4034953217;
        test_addr[2742] = 149;
        test_data[2742] = 33'd2268132089;
        test_addr[2743] = 838;
        test_data[2743] = 33'd1113939390;
        test_addr[2744] = 803;
        test_data[2744] = 33'd1913165819;
        test_addr[2745] = 746;
        test_data[2745] = 33'd2332255621;
        test_addr[2746] = 914;
        test_data[2746] = 33'd6730148341;
        test_addr[2747] = 128;
        test_data[2747] = 33'd4960252531;
        test_addr[2748] = 770;
        test_data[2748] = 33'd5198229621;
        test_addr[2749] = 424;
        test_data[2749] = 33'd6256836238;
        test_addr[2750] = 908;
        test_data[2750] = 33'd5970344877;
        test_addr[2751] = 242;
        test_data[2751] = 33'd1982815146;
        test_addr[2752] = 91;
        test_data[2752] = 33'd7566339559;
        test_addr[2753] = 1019;
        test_data[2753] = 33'd3823758254;
        test_addr[2754] = 640;
        test_data[2754] = 33'd2313811608;
        test_addr[2755] = 1023;
        test_data[2755] = 33'd6144982272;
        test_addr[2756] = 1023;
        test_data[2756] = 33'd1850014976;
        test_addr[2757] = 408;
        test_data[2757] = 33'd1130836166;
        test_addr[2758] = 20;
        test_data[2758] = 33'd4222788375;
        test_addr[2759] = 41;
        test_data[2759] = 33'd6944032070;
        test_addr[2760] = 426;
        test_data[2760] = 33'd2914022316;
        test_addr[2761] = 419;
        test_data[2761] = 33'd6344123910;
        test_addr[2762] = 196;
        test_data[2762] = 33'd1791433486;
        test_addr[2763] = 73;
        test_data[2763] = 33'd775081083;
        test_addr[2764] = 519;
        test_data[2764] = 33'd1283402259;
        test_addr[2765] = 792;
        test_data[2765] = 33'd4103913134;
        test_addr[2766] = 955;
        test_data[2766] = 33'd2326066714;
        test_addr[2767] = 846;
        test_data[2767] = 33'd7478896832;
        test_addr[2768] = 1005;
        test_data[2768] = 33'd4672360408;
        test_addr[2769] = 654;
        test_data[2769] = 33'd6910382253;
        test_addr[2770] = 713;
        test_data[2770] = 33'd333588719;
        test_addr[2771] = 211;
        test_data[2771] = 33'd3322545857;
        test_addr[2772] = 109;
        test_data[2772] = 33'd8324039898;
        test_addr[2773] = 20;
        test_data[2773] = 33'd6189677051;
        test_addr[2774] = 930;
        test_data[2774] = 33'd2007557742;
        test_addr[2775] = 93;
        test_data[2775] = 33'd6711303486;
        test_addr[2776] = 915;
        test_data[2776] = 33'd1268898235;
        test_addr[2777] = 742;
        test_data[2777] = 33'd6715008480;
        test_addr[2778] = 573;
        test_data[2778] = 33'd8195318183;
        test_addr[2779] = 433;
        test_data[2779] = 33'd5727765376;
        test_addr[2780] = 447;
        test_data[2780] = 33'd7114806516;
        test_addr[2781] = 699;
        test_data[2781] = 33'd1140078632;
        test_addr[2782] = 411;
        test_data[2782] = 33'd6426455647;
        test_addr[2783] = 811;
        test_data[2783] = 33'd712960676;
        test_addr[2784] = 434;
        test_data[2784] = 33'd188263586;
        test_addr[2785] = 1015;
        test_data[2785] = 33'd2062647632;
        test_addr[2786] = 854;
        test_data[2786] = 33'd2260897852;
        test_addr[2787] = 648;
        test_data[2787] = 33'd936482943;
        test_addr[2788] = 467;
        test_data[2788] = 33'd1242458990;
        test_addr[2789] = 196;
        test_data[2789] = 33'd5178056563;
        test_addr[2790] = 991;
        test_data[2790] = 33'd3554038044;
        test_addr[2791] = 211;
        test_data[2791] = 33'd3322545857;
        test_addr[2792] = 517;
        test_data[2792] = 33'd385111081;
        test_addr[2793] = 33;
        test_data[2793] = 33'd1484688907;
        test_addr[2794] = 569;
        test_data[2794] = 33'd2585983587;
        test_addr[2795] = 100;
        test_data[2795] = 33'd520744879;
        test_addr[2796] = 714;
        test_data[2796] = 33'd761390289;
        test_addr[2797] = 262;
        test_data[2797] = 33'd3966004824;
        test_addr[2798] = 338;
        test_data[2798] = 33'd3242582816;
        test_addr[2799] = 873;
        test_data[2799] = 33'd6159176736;
        test_addr[2800] = 558;
        test_data[2800] = 33'd4743647636;
        test_addr[2801] = 548;
        test_data[2801] = 33'd2835990504;
        test_addr[2802] = 655;
        test_data[2802] = 33'd2678884701;
        test_addr[2803] = 653;
        test_data[2803] = 33'd1819710919;
        test_addr[2804] = 565;
        test_data[2804] = 33'd7045143922;
        test_addr[2805] = 700;
        test_data[2805] = 33'd7891462331;
        test_addr[2806] = 52;
        test_data[2806] = 33'd5013461635;
        test_addr[2807] = 603;
        test_data[2807] = 33'd2447831809;
        test_addr[2808] = 506;
        test_data[2808] = 33'd3145293850;
        test_addr[2809] = 29;
        test_data[2809] = 33'd260193810;
        test_addr[2810] = 984;
        test_data[2810] = 33'd3168600535;
        test_addr[2811] = 718;
        test_data[2811] = 33'd2587264415;
        test_addr[2812] = 872;
        test_data[2812] = 33'd4939001500;
        test_addr[2813] = 729;
        test_data[2813] = 33'd1035742076;
        test_addr[2814] = 348;
        test_data[2814] = 33'd3222427471;
        test_addr[2815] = 168;
        test_data[2815] = 33'd7752897503;
        test_addr[2816] = 550;
        test_data[2816] = 33'd2861464618;
        test_addr[2817] = 479;
        test_data[2817] = 33'd6681165366;
        test_addr[2818] = 130;
        test_data[2818] = 33'd822764357;
        test_addr[2819] = 873;
        test_data[2819] = 33'd7840937683;
        test_addr[2820] = 507;
        test_data[2820] = 33'd2429522140;
        test_addr[2821] = 582;
        test_data[2821] = 33'd1527597100;
        test_addr[2822] = 803;
        test_data[2822] = 33'd1913165819;
        test_addr[2823] = 324;
        test_data[2823] = 33'd330852185;
        test_addr[2824] = 439;
        test_data[2824] = 33'd1333283651;
        test_addr[2825] = 579;
        test_data[2825] = 33'd5515249691;
        test_addr[2826] = 533;
        test_data[2826] = 33'd3809017245;
        test_addr[2827] = 587;
        test_data[2827] = 33'd702014159;
        test_addr[2828] = 410;
        test_data[2828] = 33'd3405405453;
        test_addr[2829] = 895;
        test_data[2829] = 33'd3170848996;
        test_addr[2830] = 895;
        test_data[2830] = 33'd3170848996;
        test_addr[2831] = 552;
        test_data[2831] = 33'd2630489937;
        test_addr[2832] = 546;
        test_data[2832] = 33'd555802139;
        test_addr[2833] = 638;
        test_data[2833] = 33'd8377416771;
        test_addr[2834] = 538;
        test_data[2834] = 33'd26257848;
        test_addr[2835] = 333;
        test_data[2835] = 33'd7713987545;
        test_addr[2836] = 161;
        test_data[2836] = 33'd7917722720;
        test_addr[2837] = 191;
        test_data[2837] = 33'd134572267;
        test_addr[2838] = 634;
        test_data[2838] = 33'd2731773946;
        test_addr[2839] = 318;
        test_data[2839] = 33'd1218864492;
        test_addr[2840] = 123;
        test_data[2840] = 33'd5834953353;
        test_addr[2841] = 455;
        test_data[2841] = 33'd2867352729;
        test_addr[2842] = 525;
        test_data[2842] = 33'd2628982812;
        test_addr[2843] = 665;
        test_data[2843] = 33'd1128756264;
        test_addr[2844] = 778;
        test_data[2844] = 33'd2328453822;
        test_addr[2845] = 41;
        test_data[2845] = 33'd2649064774;
        test_addr[2846] = 700;
        test_data[2846] = 33'd6868715878;
        test_addr[2847] = 261;
        test_data[2847] = 33'd2865755699;
        test_addr[2848] = 236;
        test_data[2848] = 33'd7080992697;
        test_addr[2849] = 944;
        test_data[2849] = 33'd762667074;
        test_addr[2850] = 73;
        test_data[2850] = 33'd775081083;
        test_addr[2851] = 286;
        test_data[2851] = 33'd2360048588;
        test_addr[2852] = 471;
        test_data[2852] = 33'd595140298;
        test_addr[2853] = 562;
        test_data[2853] = 33'd579089702;
        test_addr[2854] = 773;
        test_data[2854] = 33'd4379220691;
        test_addr[2855] = 719;
        test_data[2855] = 33'd8448290216;
        test_addr[2856] = 148;
        test_data[2856] = 33'd124878881;
        test_addr[2857] = 112;
        test_data[2857] = 33'd1290342635;
        test_addr[2858] = 461;
        test_data[2858] = 33'd4772081;
        test_addr[2859] = 330;
        test_data[2859] = 33'd1425051484;
        test_addr[2860] = 843;
        test_data[2860] = 33'd7679653024;
        test_addr[2861] = 971;
        test_data[2861] = 33'd634864571;
        test_addr[2862] = 143;
        test_data[2862] = 33'd6636087474;
        test_addr[2863] = 747;
        test_data[2863] = 33'd366863694;
        test_addr[2864] = 250;
        test_data[2864] = 33'd7495065624;
        test_addr[2865] = 787;
        test_data[2865] = 33'd7379110377;
        test_addr[2866] = 104;
        test_data[2866] = 33'd5650572442;
        test_addr[2867] = 729;
        test_data[2867] = 33'd1035742076;
        test_addr[2868] = 684;
        test_data[2868] = 33'd3058060985;
        test_addr[2869] = 970;
        test_data[2869] = 33'd748946215;
        test_addr[2870] = 856;
        test_data[2870] = 33'd975862316;
        test_addr[2871] = 487;
        test_data[2871] = 33'd1334951346;
        test_addr[2872] = 799;
        test_data[2872] = 33'd3954575845;
        test_addr[2873] = 28;
        test_data[2873] = 33'd8497319778;
        test_addr[2874] = 950;
        test_data[2874] = 33'd8422230215;
        test_addr[2875] = 543;
        test_data[2875] = 33'd3369326361;
        test_addr[2876] = 535;
        test_data[2876] = 33'd1384824159;
        test_addr[2877] = 145;
        test_data[2877] = 33'd1214215057;
        test_addr[2878] = 410;
        test_data[2878] = 33'd3405405453;
        test_addr[2879] = 322;
        test_data[2879] = 33'd3243207308;
        test_addr[2880] = 41;
        test_data[2880] = 33'd2649064774;
        test_addr[2881] = 407;
        test_data[2881] = 33'd1117760925;
        test_addr[2882] = 122;
        test_data[2882] = 33'd1522076612;
        test_addr[2883] = 114;
        test_data[2883] = 33'd486022466;
        test_addr[2884] = 217;
        test_data[2884] = 33'd3904384728;
        test_addr[2885] = 205;
        test_data[2885] = 33'd1920400090;
        test_addr[2886] = 166;
        test_data[2886] = 33'd1217876369;
        test_addr[2887] = 476;
        test_data[2887] = 33'd3848503637;
        test_addr[2888] = 736;
        test_data[2888] = 33'd7209479372;
        test_addr[2889] = 201;
        test_data[2889] = 33'd7021461195;
        test_addr[2890] = 266;
        test_data[2890] = 33'd8053278914;
        test_addr[2891] = 951;
        test_data[2891] = 33'd7733637949;
        test_addr[2892] = 856;
        test_data[2892] = 33'd975862316;
        test_addr[2893] = 870;
        test_data[2893] = 33'd8055043496;
        test_addr[2894] = 760;
        test_data[2894] = 33'd4199067864;
        test_addr[2895] = 733;
        test_data[2895] = 33'd3919399191;
        test_addr[2896] = 50;
        test_data[2896] = 33'd7247413534;
        test_addr[2897] = 533;
        test_data[2897] = 33'd3809017245;
        test_addr[2898] = 909;
        test_data[2898] = 33'd4376411868;
        test_addr[2899] = 278;
        test_data[2899] = 33'd3853850877;
        test_addr[2900] = 496;
        test_data[2900] = 33'd482673616;
        test_addr[2901] = 38;
        test_data[2901] = 33'd8439370794;
        test_addr[2902] = 947;
        test_data[2902] = 33'd422133090;
        test_addr[2903] = 856;
        test_data[2903] = 33'd975862316;
        test_addr[2904] = 908;
        test_data[2904] = 33'd4453686008;
        test_addr[2905] = 907;
        test_data[2905] = 33'd6471059900;
        test_addr[2906] = 412;
        test_data[2906] = 33'd1687805123;
        test_addr[2907] = 442;
        test_data[2907] = 33'd6229218759;
        test_addr[2908] = 865;
        test_data[2908] = 33'd2502908565;
        test_addr[2909] = 384;
        test_data[2909] = 33'd2775621126;
        test_addr[2910] = 708;
        test_data[2910] = 33'd3363550927;
        test_addr[2911] = 433;
        test_data[2911] = 33'd1432798080;
        test_addr[2912] = 850;
        test_data[2912] = 33'd640217809;
        test_addr[2913] = 283;
        test_data[2913] = 33'd581010001;
        test_addr[2914] = 40;
        test_data[2914] = 33'd2224301287;
        test_addr[2915] = 791;
        test_data[2915] = 33'd1738721985;
        test_addr[2916] = 64;
        test_data[2916] = 33'd3038722049;
        test_addr[2917] = 1009;
        test_data[2917] = 33'd4723747292;
        test_addr[2918] = 694;
        test_data[2918] = 33'd620562415;
        test_addr[2919] = 199;
        test_data[2919] = 33'd8483066573;
        test_addr[2920] = 771;
        test_data[2920] = 33'd5053070985;
        test_addr[2921] = 87;
        test_data[2921] = 33'd6670938754;
        test_addr[2922] = 818;
        test_data[2922] = 33'd4648027946;
        test_addr[2923] = 324;
        test_data[2923] = 33'd6071292160;
        test_addr[2924] = 76;
        test_data[2924] = 33'd3779515059;
        test_addr[2925] = 695;
        test_data[2925] = 33'd2186911345;
        test_addr[2926] = 1017;
        test_data[2926] = 33'd7592464259;
        test_addr[2927] = 193;
        test_data[2927] = 33'd8054981974;
        test_addr[2928] = 723;
        test_data[2928] = 33'd5020869985;
        test_addr[2929] = 146;
        test_data[2929] = 33'd3440025518;
        test_addr[2930] = 977;
        test_data[2930] = 33'd5188510135;
        test_addr[2931] = 510;
        test_data[2931] = 33'd363583401;
        test_addr[2932] = 682;
        test_data[2932] = 33'd301906037;
        test_addr[2933] = 242;
        test_data[2933] = 33'd7749610354;
        test_addr[2934] = 588;
        test_data[2934] = 33'd4041263385;
        test_addr[2935] = 922;
        test_data[2935] = 33'd715587172;
        test_addr[2936] = 1016;
        test_data[2936] = 33'd1926784674;
        test_addr[2937] = 89;
        test_data[2937] = 33'd201002197;
        test_addr[2938] = 539;
        test_data[2938] = 33'd3811829804;
        test_addr[2939] = 519;
        test_data[2939] = 33'd7767383272;
        test_addr[2940] = 858;
        test_data[2940] = 33'd1025625720;
        test_addr[2941] = 165;
        test_data[2941] = 33'd5509706080;
        test_addr[2942] = 617;
        test_data[2942] = 33'd7924547456;
        test_addr[2943] = 676;
        test_data[2943] = 33'd1174454579;
        test_addr[2944] = 194;
        test_data[2944] = 33'd2912051046;
        test_addr[2945] = 908;
        test_data[2945] = 33'd158718712;
        test_addr[2946] = 91;
        test_data[2946] = 33'd3271372263;
        test_addr[2947] = 589;
        test_data[2947] = 33'd7395626761;
        test_addr[2948] = 384;
        test_data[2948] = 33'd2775621126;
        test_addr[2949] = 693;
        test_data[2949] = 33'd2069998988;
        test_addr[2950] = 926;
        test_data[2950] = 33'd3522717221;
        test_addr[2951] = 183;
        test_data[2951] = 33'd3711706094;
        test_addr[2952] = 792;
        test_data[2952] = 33'd5266502348;
        test_addr[2953] = 619;
        test_data[2953] = 33'd5653505965;
        test_addr[2954] = 980;
        test_data[2954] = 33'd8193866474;
        test_addr[2955] = 318;
        test_data[2955] = 33'd1218864492;
        test_addr[2956] = 759;
        test_data[2956] = 33'd2196879887;
        test_addr[2957] = 677;
        test_data[2957] = 33'd2985165387;
        test_addr[2958] = 323;
        test_data[2958] = 33'd1032448390;
        test_addr[2959] = 322;
        test_data[2959] = 33'd3243207308;
        test_addr[2960] = 538;
        test_data[2960] = 33'd26257848;
        test_addr[2961] = 871;
        test_data[2961] = 33'd7749521884;
        test_addr[2962] = 549;
        test_data[2962] = 33'd1304665201;
        test_addr[2963] = 242;
        test_data[2963] = 33'd3454643058;
        test_addr[2964] = 543;
        test_data[2964] = 33'd3369326361;
        test_addr[2965] = 118;
        test_data[2965] = 33'd4130850739;
        test_addr[2966] = 484;
        test_data[2966] = 33'd8299586646;
        test_addr[2967] = 456;
        test_data[2967] = 33'd4701616139;
        test_addr[2968] = 491;
        test_data[2968] = 33'd3769941878;
        test_addr[2969] = 781;
        test_data[2969] = 33'd8463092087;
        test_addr[2970] = 100;
        test_data[2970] = 33'd520744879;
        test_addr[2971] = 310;
        test_data[2971] = 33'd3692301779;
        test_addr[2972] = 152;
        test_data[2972] = 33'd4105911548;
        test_addr[2973] = 871;
        test_data[2973] = 33'd3454554588;
        test_addr[2974] = 322;
        test_data[2974] = 33'd3243207308;
        test_addr[2975] = 1009;
        test_data[2975] = 33'd5859866907;
        test_addr[2976] = 958;
        test_data[2976] = 33'd3257284543;
        test_addr[2977] = 35;
        test_data[2977] = 33'd2325257392;
        test_addr[2978] = 505;
        test_data[2978] = 33'd6546109174;
        test_addr[2979] = 793;
        test_data[2979] = 33'd1650429696;
        test_addr[2980] = 973;
        test_data[2980] = 33'd986805218;
        test_addr[2981] = 25;
        test_data[2981] = 33'd2605255280;
        test_addr[2982] = 298;
        test_data[2982] = 33'd1530159267;
        test_addr[2983] = 248;
        test_data[2983] = 33'd6868030587;
        test_addr[2984] = 900;
        test_data[2984] = 33'd3715729542;
        test_addr[2985] = 105;
        test_data[2985] = 33'd3407001355;
        test_addr[2986] = 132;
        test_data[2986] = 33'd5559059375;
        test_addr[2987] = 174;
        test_data[2987] = 33'd3604100316;
        test_addr[2988] = 153;
        test_data[2988] = 33'd632865373;
        test_addr[2989] = 505;
        test_data[2989] = 33'd5326281240;
        test_addr[2990] = 412;
        test_data[2990] = 33'd8541409316;
        test_addr[2991] = 140;
        test_data[2991] = 33'd3162183515;
        test_addr[2992] = 618;
        test_data[2992] = 33'd5461278113;
        test_addr[2993] = 285;
        test_data[2993] = 33'd1566790510;
        test_addr[2994] = 139;
        test_data[2994] = 33'd4181971414;
        test_addr[2995] = 561;
        test_data[2995] = 33'd1350524622;
        test_addr[2996] = 979;
        test_data[2996] = 33'd7755950886;
        test_addr[2997] = 386;
        test_data[2997] = 33'd1131231838;
        test_addr[2998] = 738;
        test_data[2998] = 33'd841875993;
        test_addr[2999] = 681;
        test_data[2999] = 33'd1711100772;

    end
endmodule


/*
本文件是一个测试文件，用于测试cache模块
工作原理是模仿CPU的读写请求，对cache进行读写操作
将Cache返回的数据与预先数据进行比较，如果一致则测试通过
*/
`timescale 1ns/1ps
module cache_tb();

    //测试参数
    parameter READ_NUM = 2000;  // 测试次数 这里设置为2000次读，1000次写
    parameter WRITE_NUM = 1000;  
    //模块参数
    parameter INDEX_WIDTH       = 3;   // Cache索引位宽 2^3=8行
    parameter LINE_OFFSET_WIDTH = 2;   // 行偏移位宽，决定了一行的宽度 2^2=4字
    parameter SPACE_OFFSET      = 2;   // 一个地址空间占1个字节，因此一个字需要4个地址空间，由于假设为整字读取，处理地址的时候可以默认后两位为0
    parameter MEM_ADDR_WIDTH    = 10;   // 为了简化，这里假设内存地址宽度为10位（CPU请求地址仍然是32位，只不过我们这里简化处理，截断了高位） 
    parameter WAY_NUM           = 2;   // Cache N路组相联(N=1的时候是直接映射)
    parameter REPLACE_POLICY    = 0;   // 替换策略 0：LRU 1：FIFO 2：伪随机

    // 变化的信号 CPU发出
    reg clk=1;
    reg rstn=1;
    reg stat=0;
    // 等rstn信号稳定后 clk信号才开始翻转
    initial begin
        #1 rstn = 0;
        #1 rstn = 1;
        stat = 1;
    end
    always  #1 clk = ~clk;

    wire [31:0] addr;
    wire r_req;
    wire w_req;
    wire [31:0] w_data;

    // 导线
    wire [31:0] r_data;
    wire miss;
    wire mem_r;
    wire mem_w;
    wire [31:0] mem_addr;
    wire [127:0] mem_w_data;
    wire [127:0] mem_r_data;
    wire mem_ready;

    // 用于测试的信号
    reg [MEM_ADDR_WIDTH-1:0] test_addr[0:READ_NUM+WRITE_NUM-1];  // 用于存储测试地址
    reg [32:0] test_data[0:READ_NUM+WRITE_NUM-1];  // 用于存储测试数据 最高位用于标记是否写入 0：读 1：写
    reg [31:0] test_cnt=0;  // 用于计数，每次读写操作后加1
    reg diff=0;  // 用于标记是否有不一致的数据

    // 用于对比的提交，当前cache应该给出的数据
    wire op;
    wire[31:0] data;
    assign op = test_data[test_cnt-1][32];
    assign data = test_data[test_cnt-1][31:0];
    
    // 状态机
    assign addr = test_addr[test_cnt]<<SPACE_OFFSET;
    assign r_req = test_data[test_cnt][32] == 0 ? 1 : 0;
    assign w_req = test_data[test_cnt][32] == 1 ? 1 : 0;
    assign w_data = test_data[test_cnt][31:0];
    always @(posedge clk) begin
        if (!miss && (test_cnt < READ_NUM+WRITE_NUM) && stat) begin
            if (test_data[test_cnt-1][32] == 0) begin  // 读
                if (r_data != test_data[test_cnt-1][31:0]) begin
                    $display("Read error at %d, expect %h, get %h", test_cnt, test_data[test_cnt-1][31:0], r_data);
                    diff = 1;
                end
            end
            test_cnt <= test_cnt + 1;
        end
    end

    // 例化cache
    cache #(
        .INDEX_WIDTH(INDEX_WIDTH),
        .LINE_OFFSET_WIDTH(LINE_OFFSET_WIDTH),
        .SPACE_OFFSET(SPACE_OFFSET),
        .WAY_NUM(WAY_NUM),
        .REPLACE_POLICY(REPLACE_POLICY)
    ) cache_inst(
        .clk(clk),
        .rstn(rstn),
        .addr(addr),
        .r_req(r_req),
        .w_req(w_req),
        .w_data(w_data),
        .r_data(r_data),
        .miss(miss),
        .mem_r(mem_r),
        .mem_w(mem_w),
        .mem_addr(mem_addr),
        .mem_w_data(mem_w_data),
        .mem_r_data(mem_r_data),
        .mem_ready(mem_ready)
    );

    // 内存
    mem #(
        .INDEX_WIDTH(INDEX_WIDTH),
        .LINE_OFFSET_WIDTH(LINE_OFFSET_WIDTH),
        .SPACE_OFFSET(SPACE_OFFSET),
        .MEM_ADDR_WIDTH(MEM_ADDR_WIDTH-LINE_OFFSET_WIDTH),
        .WAY_NUM(WAY_NUM)
    ) mem_inst(
        .clk(clk),
        .rstn(rstn),
        .mem_r(mem_r),
        .mem_w(mem_w),
        .mem_addr(mem_addr),
        .mem_w_data(mem_w_data),
        .mem_r_data(mem_r_data),
        .mem_ready(mem_ready)
    );

    // 初始化测试数据
    initial begin
        test_addr[0] = 0;
        test_data[0] = 33'd1870585436;
        test_addr[1] = 1;
        test_data[1] = 33'd6159452856;
        test_addr[2] = 2;
        test_data[2] = 33'd6248579081;
        test_addr[3] = 3;
        test_data[3] = 33'd3350406635;
        test_addr[4] = 4;
        test_data[4] = 33'd5758728835;
        test_addr[5] = 5;
        test_data[5] = 33'd2154190107;
        test_addr[6] = 6;
        test_data[6] = 33'd5889149421;
        test_addr[7] = 7;
        test_data[7] = 33'd4633379770;
        test_addr[8] = 8;
        test_data[8] = 33'd3505230681;
        test_addr[9] = 9;
        test_data[9] = 33'd5667747975;
        test_addr[10] = 606;
        test_data[10] = 33'd906696308;
        test_addr[11] = 607;
        test_data[11] = 33'd7980303264;
        test_addr[12] = 608;
        test_data[12] = 33'd3635138265;
        test_addr[13] = 10;
        test_data[13] = 33'd4271687727;
        test_addr[14] = 11;
        test_data[14] = 33'd2298463057;
        test_addr[15] = 309;
        test_data[15] = 33'd3941608837;
        test_addr[16] = 310;
        test_data[16] = 33'd3094631771;
        test_addr[17] = 311;
        test_data[17] = 33'd1449524691;
        test_addr[18] = 312;
        test_data[18] = 33'd240548675;
        test_addr[19] = 313;
        test_data[19] = 33'd7364133990;
        test_addr[20] = 314;
        test_data[20] = 33'd3194236288;
        test_addr[21] = 315;
        test_data[21] = 33'd3309303920;
        test_addr[22] = 316;
        test_data[22] = 33'd838957123;
        test_addr[23] = 317;
        test_data[23] = 33'd8407323568;
        test_addr[24] = 318;
        test_data[24] = 33'd5662154682;
        test_addr[25] = 319;
        test_data[25] = 33'd4693333721;
        test_addr[26] = 320;
        test_data[26] = 33'd6508072877;
        test_addr[27] = 321;
        test_data[27] = 33'd4078285937;
        test_addr[28] = 322;
        test_data[28] = 33'd4172724571;
        test_addr[29] = 323;
        test_data[29] = 33'd2407757486;
        test_addr[30] = 324;
        test_data[30] = 33'd6734438521;
        test_addr[31] = 325;
        test_data[31] = 33'd7290604514;
        test_addr[32] = 326;
        test_data[32] = 33'd7326668415;
        test_addr[33] = 327;
        test_data[33] = 33'd318989378;
        test_addr[34] = 328;
        test_data[34] = 33'd3131202390;
        test_addr[35] = 329;
        test_data[35] = 33'd5732614156;
        test_addr[36] = 330;
        test_data[36] = 33'd1703867803;
        test_addr[37] = 331;
        test_data[37] = 33'd2887064224;
        test_addr[38] = 332;
        test_data[38] = 33'd3238606923;
        test_addr[39] = 333;
        test_data[39] = 33'd5757291551;
        test_addr[40] = 334;
        test_data[40] = 33'd8204252092;
        test_addr[41] = 12;
        test_data[41] = 33'd1768449257;
        test_addr[42] = 13;
        test_data[42] = 33'd4162140124;
        test_addr[43] = 14;
        test_data[43] = 33'd539032534;
        test_addr[44] = 15;
        test_data[44] = 33'd1119003857;
        test_addr[45] = 16;
        test_data[45] = 33'd3925987810;
        test_addr[46] = 17;
        test_data[46] = 33'd1949417226;
        test_addr[47] = 18;
        test_data[47] = 33'd1569000094;
        test_addr[48] = 19;
        test_data[48] = 33'd7618478519;
        test_addr[49] = 20;
        test_data[49] = 33'd592586045;
        test_addr[50] = 21;
        test_data[50] = 33'd5496505057;
        test_addr[51] = 22;
        test_data[51] = 33'd1621961986;
        test_addr[52] = 23;
        test_data[52] = 33'd4536436496;
        test_addr[53] = 24;
        test_data[53] = 33'd2159349817;
        test_addr[54] = 25;
        test_data[54] = 33'd7768116034;
        test_addr[55] = 26;
        test_data[55] = 33'd7317503360;
        test_addr[56] = 27;
        test_data[56] = 33'd1798709310;
        test_addr[57] = 28;
        test_data[57] = 33'd4030679079;
        test_addr[58] = 29;
        test_data[58] = 33'd3629881189;
        test_addr[59] = 30;
        test_data[59] = 33'd1193996624;
        test_addr[60] = 31;
        test_data[60] = 33'd3527005491;
        test_addr[61] = 32;
        test_data[61] = 33'd3844512050;
        test_addr[62] = 33;
        test_data[62] = 33'd6718771741;
        test_addr[63] = 34;
        test_data[63] = 33'd1289644746;
        test_addr[64] = 35;
        test_data[64] = 33'd1604560142;
        test_addr[65] = 36;
        test_data[65] = 33'd5736960618;
        test_addr[66] = 37;
        test_data[66] = 33'd3077452828;
        test_addr[67] = 38;
        test_data[67] = 33'd179744430;
        test_addr[68] = 39;
        test_data[68] = 33'd8569920432;
        test_addr[69] = 40;
        test_data[69] = 33'd1444412845;
        test_addr[70] = 41;
        test_data[70] = 33'd660859156;
        test_addr[71] = 42;
        test_data[71] = 33'd6562869273;
        test_addr[72] = 43;
        test_data[72] = 33'd5893661504;
        test_addr[73] = 44;
        test_data[73] = 33'd4793613235;
        test_addr[74] = 45;
        test_data[74] = 33'd7052709041;
        test_addr[75] = 46;
        test_data[75] = 33'd4612300498;
        test_addr[76] = 47;
        test_data[76] = 33'd999277383;
        test_addr[77] = 45;
        test_data[77] = 33'd2757741745;
        test_addr[78] = 46;
        test_data[78] = 33'd317333202;
        test_addr[79] = 47;
        test_data[79] = 33'd999277383;
        test_addr[80] = 48;
        test_data[80] = 33'd2577690104;
        test_addr[81] = 49;
        test_data[81] = 33'd2828154457;
        test_addr[82] = 50;
        test_data[82] = 33'd3713624851;
        test_addr[83] = 51;
        test_data[83] = 33'd3352351002;
        test_addr[84] = 52;
        test_data[84] = 33'd3291818831;
        test_addr[85] = 53;
        test_data[85] = 33'd48823010;
        test_addr[86] = 54;
        test_data[86] = 33'd1614540136;
        test_addr[87] = 55;
        test_data[87] = 33'd4041042842;
        test_addr[88] = 56;
        test_data[88] = 33'd2473651066;
        test_addr[89] = 57;
        test_data[89] = 33'd400692079;
        test_addr[90] = 58;
        test_data[90] = 33'd2831688436;
        test_addr[91] = 59;
        test_data[91] = 33'd1487397129;
        test_addr[92] = 60;
        test_data[92] = 33'd6381573462;
        test_addr[93] = 61;
        test_data[93] = 33'd3519769342;
        test_addr[94] = 62;
        test_data[94] = 33'd504570280;
        test_addr[95] = 63;
        test_data[95] = 33'd2384061833;
        test_addr[96] = 64;
        test_data[96] = 33'd4168218661;
        test_addr[97] = 65;
        test_data[97] = 33'd8464452811;
        test_addr[98] = 66;
        test_data[98] = 33'd876819121;
        test_addr[99] = 48;
        test_data[99] = 33'd2577690104;
        test_addr[100] = 49;
        test_data[100] = 33'd7176035497;
        test_addr[101] = 50;
        test_data[101] = 33'd6612078940;
        test_addr[102] = 51;
        test_data[102] = 33'd3352351002;
        test_addr[103] = 52;
        test_data[103] = 33'd3291818831;
        test_addr[104] = 53;
        test_data[104] = 33'd48823010;
        test_addr[105] = 54;
        test_data[105] = 33'd1614540136;
        test_addr[106] = 55;
        test_data[106] = 33'd8488122069;
        test_addr[107] = 56;
        test_data[107] = 33'd2473651066;
        test_addr[108] = 57;
        test_data[108] = 33'd4316978358;
        test_addr[109] = 58;
        test_data[109] = 33'd7498115080;
        test_addr[110] = 59;
        test_data[110] = 33'd1487397129;
        test_addr[111] = 60;
        test_data[111] = 33'd2086606166;
        test_addr[112] = 741;
        test_data[112] = 33'd1810153704;
        test_addr[113] = 742;
        test_data[113] = 33'd2878401245;
        test_addr[114] = 743;
        test_data[114] = 33'd292010483;
        test_addr[115] = 744;
        test_data[115] = 33'd230455895;
        test_addr[116] = 745;
        test_data[116] = 33'd3435630877;
        test_addr[117] = 746;
        test_data[117] = 33'd3185922216;
        test_addr[118] = 747;
        test_data[118] = 33'd7744800262;
        test_addr[119] = 748;
        test_data[119] = 33'd3916469345;
        test_addr[120] = 749;
        test_data[120] = 33'd1248251572;
        test_addr[121] = 61;
        test_data[121] = 33'd6830345116;
        test_addr[122] = 62;
        test_data[122] = 33'd504570280;
        test_addr[123] = 63;
        test_data[123] = 33'd2384061833;
        test_addr[124] = 64;
        test_data[124] = 33'd4168218661;
        test_addr[125] = 65;
        test_data[125] = 33'd4169485515;
        test_addr[126] = 66;
        test_data[126] = 33'd876819121;
        test_addr[127] = 67;
        test_data[127] = 33'd2886172558;
        test_addr[128] = 68;
        test_data[128] = 33'd6735359636;
        test_addr[129] = 69;
        test_data[129] = 33'd5007320758;
        test_addr[130] = 70;
        test_data[130] = 33'd3874690545;
        test_addr[131] = 71;
        test_data[131] = 33'd6095592192;
        test_addr[132] = 72;
        test_data[132] = 33'd8040442258;
        test_addr[133] = 73;
        test_data[133] = 33'd6770459619;
        test_addr[134] = 74;
        test_data[134] = 33'd3146623705;
        test_addr[135] = 75;
        test_data[135] = 33'd3972422453;
        test_addr[136] = 76;
        test_data[136] = 33'd1051232611;
        test_addr[137] = 77;
        test_data[137] = 33'd998193764;
        test_addr[138] = 78;
        test_data[138] = 33'd3095344887;
        test_addr[139] = 79;
        test_data[139] = 33'd466432104;
        test_addr[140] = 80;
        test_data[140] = 33'd3440150321;
        test_addr[141] = 81;
        test_data[141] = 33'd2716768050;
        test_addr[142] = 82;
        test_data[142] = 33'd979668869;
        test_addr[143] = 83;
        test_data[143] = 33'd7767129141;
        test_addr[144] = 84;
        test_data[144] = 33'd4684736685;
        test_addr[145] = 491;
        test_data[145] = 33'd8565251703;
        test_addr[146] = 85;
        test_data[146] = 33'd3703089126;
        test_addr[147] = 86;
        test_data[147] = 33'd623629618;
        test_addr[148] = 69;
        test_data[148] = 33'd712353462;
        test_addr[149] = 70;
        test_data[149] = 33'd3874690545;
        test_addr[150] = 71;
        test_data[150] = 33'd1800624896;
        test_addr[151] = 72;
        test_data[151] = 33'd3745474962;
        test_addr[152] = 73;
        test_data[152] = 33'd7885172759;
        test_addr[153] = 74;
        test_data[153] = 33'd3146623705;
        test_addr[154] = 75;
        test_data[154] = 33'd3972422453;
        test_addr[155] = 76;
        test_data[155] = 33'd1051232611;
        test_addr[156] = 77;
        test_data[156] = 33'd998193764;
        test_addr[157] = 78;
        test_data[157] = 33'd7886457610;
        test_addr[158] = 79;
        test_data[158] = 33'd466432104;
        test_addr[159] = 80;
        test_data[159] = 33'd3440150321;
        test_addr[160] = 81;
        test_data[160] = 33'd6904617404;
        test_addr[161] = 82;
        test_data[161] = 33'd5027633604;
        test_addr[162] = 83;
        test_data[162] = 33'd3472161845;
        test_addr[163] = 84;
        test_data[163] = 33'd389769389;
        test_addr[164] = 87;
        test_data[164] = 33'd3303907992;
        test_addr[165] = 88;
        test_data[165] = 33'd1506464650;
        test_addr[166] = 89;
        test_data[166] = 33'd1036241526;
        test_addr[167] = 90;
        test_data[167] = 33'd548807498;
        test_addr[168] = 91;
        test_data[168] = 33'd3415150818;
        test_addr[169] = 92;
        test_data[169] = 33'd4105109197;
        test_addr[170] = 93;
        test_data[170] = 33'd4048368480;
        test_addr[171] = 94;
        test_data[171] = 33'd2640578934;
        test_addr[172] = 95;
        test_data[172] = 33'd6518326159;
        test_addr[173] = 96;
        test_data[173] = 33'd1607774016;
        test_addr[174] = 97;
        test_data[174] = 33'd2681259618;
        test_addr[175] = 98;
        test_data[175] = 33'd1885671812;
        test_addr[176] = 99;
        test_data[176] = 33'd2668054470;
        test_addr[177] = 100;
        test_data[177] = 33'd3329548407;
        test_addr[178] = 101;
        test_data[178] = 33'd5825670757;
        test_addr[179] = 102;
        test_data[179] = 33'd7927049670;
        test_addr[180] = 103;
        test_data[180] = 33'd7202537296;
        test_addr[181] = 104;
        test_data[181] = 33'd6699030592;
        test_addr[182] = 331;
        test_data[182] = 33'd2887064224;
        test_addr[183] = 332;
        test_data[183] = 33'd3238606923;
        test_addr[184] = 333;
        test_data[184] = 33'd1462324255;
        test_addr[185] = 334;
        test_data[185] = 33'd3909284796;
        test_addr[186] = 335;
        test_data[186] = 33'd115410482;
        test_addr[187] = 336;
        test_data[187] = 33'd2188727585;
        test_addr[188] = 337;
        test_data[188] = 33'd325795203;
        test_addr[189] = 338;
        test_data[189] = 33'd3556465203;
        test_addr[190] = 339;
        test_data[190] = 33'd2720908177;
        test_addr[191] = 340;
        test_data[191] = 33'd5925762037;
        test_addr[192] = 341;
        test_data[192] = 33'd829190514;
        test_addr[193] = 342;
        test_data[193] = 33'd2723057950;
        test_addr[194] = 343;
        test_data[194] = 33'd5931483359;
        test_addr[195] = 344;
        test_data[195] = 33'd281373290;
        test_addr[196] = 345;
        test_data[196] = 33'd3249490296;
        test_addr[197] = 346;
        test_data[197] = 33'd3397465739;
        test_addr[198] = 347;
        test_data[198] = 33'd184952467;
        test_addr[199] = 348;
        test_data[199] = 33'd7396581503;
        test_addr[200] = 349;
        test_data[200] = 33'd4811787517;
        test_addr[201] = 350;
        test_data[201] = 33'd5413869609;
        test_addr[202] = 351;
        test_data[202] = 33'd5212194063;
        test_addr[203] = 352;
        test_data[203] = 33'd147931898;
        test_addr[204] = 353;
        test_data[204] = 33'd1647595599;
        test_addr[205] = 354;
        test_data[205] = 33'd3966319412;
        test_addr[206] = 355;
        test_data[206] = 33'd7569737053;
        test_addr[207] = 356;
        test_data[207] = 33'd3033278383;
        test_addr[208] = 357;
        test_data[208] = 33'd5394600868;
        test_addr[209] = 358;
        test_data[209] = 33'd928067253;
        test_addr[210] = 359;
        test_data[210] = 33'd4082684122;
        test_addr[211] = 360;
        test_data[211] = 33'd1883443685;
        test_addr[212] = 361;
        test_data[212] = 33'd5146389209;
        test_addr[213] = 362;
        test_data[213] = 33'd3612932426;
        test_addr[214] = 363;
        test_data[214] = 33'd3770020475;
        test_addr[215] = 364;
        test_data[215] = 33'd4047546126;
        test_addr[216] = 365;
        test_data[216] = 33'd4577362485;
        test_addr[217] = 366;
        test_data[217] = 33'd2115114658;
        test_addr[218] = 367;
        test_data[218] = 33'd5211361410;
        test_addr[219] = 368;
        test_data[219] = 33'd3673022184;
        test_addr[220] = 369;
        test_data[220] = 33'd4682027180;
        test_addr[221] = 370;
        test_data[221] = 33'd7122206462;
        test_addr[222] = 371;
        test_data[222] = 33'd4593873379;
        test_addr[223] = 105;
        test_data[223] = 33'd1914703890;
        test_addr[224] = 501;
        test_data[224] = 33'd2750530624;
        test_addr[225] = 502;
        test_data[225] = 33'd6724105452;
        test_addr[226] = 503;
        test_data[226] = 33'd5445741866;
        test_addr[227] = 504;
        test_data[227] = 33'd5245995105;
        test_addr[228] = 505;
        test_data[228] = 33'd1706057765;
        test_addr[229] = 506;
        test_data[229] = 33'd846958545;
        test_addr[230] = 507;
        test_data[230] = 33'd640223175;
        test_addr[231] = 508;
        test_data[231] = 33'd8074643234;
        test_addr[232] = 509;
        test_data[232] = 33'd5543024920;
        test_addr[233] = 510;
        test_data[233] = 33'd154773377;
        test_addr[234] = 511;
        test_data[234] = 33'd7637937715;
        test_addr[235] = 512;
        test_data[235] = 33'd283576485;
        test_addr[236] = 513;
        test_data[236] = 33'd3832833658;
        test_addr[237] = 514;
        test_data[237] = 33'd1019661124;
        test_addr[238] = 515;
        test_data[238] = 33'd4175963926;
        test_addr[239] = 516;
        test_data[239] = 33'd2970200192;
        test_addr[240] = 517;
        test_data[240] = 33'd5468332933;
        test_addr[241] = 518;
        test_data[241] = 33'd6719558744;
        test_addr[242] = 519;
        test_data[242] = 33'd6767028449;
        test_addr[243] = 520;
        test_data[243] = 33'd2499178703;
        test_addr[244] = 106;
        test_data[244] = 33'd4863713336;
        test_addr[245] = 619;
        test_data[245] = 33'd2051461989;
        test_addr[246] = 620;
        test_data[246] = 33'd3343656720;
        test_addr[247] = 621;
        test_data[247] = 33'd723470077;
        test_addr[248] = 107;
        test_data[248] = 33'd2329785644;
        test_addr[249] = 108;
        test_data[249] = 33'd7428887775;
        test_addr[250] = 109;
        test_data[250] = 33'd2828290416;
        test_addr[251] = 110;
        test_data[251] = 33'd7913982309;
        test_addr[252] = 839;
        test_data[252] = 33'd1323733114;
        test_addr[253] = 840;
        test_data[253] = 33'd4757912404;
        test_addr[254] = 841;
        test_data[254] = 33'd729735648;
        test_addr[255] = 842;
        test_data[255] = 33'd3905935845;
        test_addr[256] = 843;
        test_data[256] = 33'd64812169;
        test_addr[257] = 844;
        test_data[257] = 33'd1905889562;
        test_addr[258] = 845;
        test_data[258] = 33'd7219442558;
        test_addr[259] = 846;
        test_data[259] = 33'd3157279990;
        test_addr[260] = 847;
        test_data[260] = 33'd4178636307;
        test_addr[261] = 848;
        test_data[261] = 33'd1091101872;
        test_addr[262] = 849;
        test_data[262] = 33'd2875037109;
        test_addr[263] = 850;
        test_data[263] = 33'd1086596891;
        test_addr[264] = 851;
        test_data[264] = 33'd30109657;
        test_addr[265] = 852;
        test_data[265] = 33'd201249939;
        test_addr[266] = 853;
        test_data[266] = 33'd5077809495;
        test_addr[267] = 111;
        test_data[267] = 33'd2224133112;
        test_addr[268] = 269;
        test_data[268] = 33'd3243925981;
        test_addr[269] = 112;
        test_data[269] = 33'd5906202983;
        test_addr[270] = 113;
        test_data[270] = 33'd2509755899;
        test_addr[271] = 114;
        test_data[271] = 33'd759874881;
        test_addr[272] = 115;
        test_data[272] = 33'd1862517686;
        test_addr[273] = 116;
        test_data[273] = 33'd1148833960;
        test_addr[274] = 117;
        test_data[274] = 33'd1057530362;
        test_addr[275] = 118;
        test_data[275] = 33'd2857138427;
        test_addr[276] = 119;
        test_data[276] = 33'd2989373656;
        test_addr[277] = 120;
        test_data[277] = 33'd132670189;
        test_addr[278] = 121;
        test_data[278] = 33'd371426538;
        test_addr[279] = 122;
        test_data[279] = 33'd1367201542;
        test_addr[280] = 123;
        test_data[280] = 33'd4608826659;
        test_addr[281] = 124;
        test_data[281] = 33'd1496960271;
        test_addr[282] = 125;
        test_data[282] = 33'd1825838587;
        test_addr[283] = 126;
        test_data[283] = 33'd4895627930;
        test_addr[284] = 127;
        test_data[284] = 33'd415964961;
        test_addr[285] = 128;
        test_data[285] = 33'd6956675663;
        test_addr[286] = 129;
        test_data[286] = 33'd1885285401;
        test_addr[287] = 130;
        test_data[287] = 33'd454112648;
        test_addr[288] = 131;
        test_data[288] = 33'd351680695;
        test_addr[289] = 132;
        test_data[289] = 33'd4027336748;
        test_addr[290] = 133;
        test_data[290] = 33'd1549772363;
        test_addr[291] = 134;
        test_data[291] = 33'd4695543826;
        test_addr[292] = 135;
        test_data[292] = 33'd1960021159;
        test_addr[293] = 136;
        test_data[293] = 33'd3552771192;
        test_addr[294] = 137;
        test_data[294] = 33'd3115074711;
        test_addr[295] = 138;
        test_data[295] = 33'd2291202182;
        test_addr[296] = 8;
        test_data[296] = 33'd6037753470;
        test_addr[297] = 9;
        test_data[297] = 33'd8558680781;
        test_addr[298] = 10;
        test_data[298] = 33'd4271687727;
        test_addr[299] = 11;
        test_data[299] = 33'd8262722102;
        test_addr[300] = 12;
        test_data[300] = 33'd1768449257;
        test_addr[301] = 13;
        test_data[301] = 33'd5011439423;
        test_addr[302] = 14;
        test_data[302] = 33'd539032534;
        test_addr[303] = 15;
        test_data[303] = 33'd1119003857;
        test_addr[304] = 16;
        test_data[304] = 33'd3925987810;
        test_addr[305] = 17;
        test_data[305] = 33'd5575695920;
        test_addr[306] = 18;
        test_data[306] = 33'd1569000094;
        test_addr[307] = 19;
        test_data[307] = 33'd3323511223;
        test_addr[308] = 20;
        test_data[308] = 33'd4512505631;
        test_addr[309] = 139;
        test_data[309] = 33'd4938753042;
        test_addr[310] = 140;
        test_data[310] = 33'd684175502;
        test_addr[311] = 141;
        test_data[311] = 33'd3385276041;
        test_addr[312] = 142;
        test_data[312] = 33'd7184726426;
        test_addr[313] = 143;
        test_data[313] = 33'd1761678698;
        test_addr[314] = 144;
        test_data[314] = 33'd7879410931;
        test_addr[315] = 145;
        test_data[315] = 33'd2276121759;
        test_addr[316] = 146;
        test_data[316] = 33'd1978812597;
        test_addr[317] = 147;
        test_data[317] = 33'd3498313420;
        test_addr[318] = 148;
        test_data[318] = 33'd8309600936;
        test_addr[319] = 149;
        test_data[319] = 33'd7634250154;
        test_addr[320] = 150;
        test_data[320] = 33'd1729930243;
        test_addr[321] = 151;
        test_data[321] = 33'd5097020712;
        test_addr[322] = 152;
        test_data[322] = 33'd5528147243;
        test_addr[323] = 153;
        test_data[323] = 33'd352254805;
        test_addr[324] = 184;
        test_data[324] = 33'd961772350;
        test_addr[325] = 185;
        test_data[325] = 33'd6740845502;
        test_addr[326] = 186;
        test_data[326] = 33'd6470528786;
        test_addr[327] = 187;
        test_data[327] = 33'd3131077888;
        test_addr[328] = 188;
        test_data[328] = 33'd4423463387;
        test_addr[329] = 189;
        test_data[329] = 33'd133639369;
        test_addr[330] = 190;
        test_data[330] = 33'd4284820396;
        test_addr[331] = 191;
        test_data[331] = 33'd7445732373;
        test_addr[332] = 192;
        test_data[332] = 33'd6890772625;
        test_addr[333] = 193;
        test_data[333] = 33'd4758040441;
        test_addr[334] = 194;
        test_data[334] = 33'd2242595831;
        test_addr[335] = 195;
        test_data[335] = 33'd186646160;
        test_addr[336] = 196;
        test_data[336] = 33'd6106370174;
        test_addr[337] = 197;
        test_data[337] = 33'd7850347484;
        test_addr[338] = 154;
        test_data[338] = 33'd4717991679;
        test_addr[339] = 155;
        test_data[339] = 33'd979919250;
        test_addr[340] = 156;
        test_data[340] = 33'd5619788673;
        test_addr[341] = 157;
        test_data[341] = 33'd1981510702;
        test_addr[342] = 158;
        test_data[342] = 33'd2395849516;
        test_addr[343] = 159;
        test_data[343] = 33'd4008254182;
        test_addr[344] = 49;
        test_data[344] = 33'd5244150990;
        test_addr[345] = 50;
        test_data[345] = 33'd8322614327;
        test_addr[346] = 51;
        test_data[346] = 33'd3352351002;
        test_addr[347] = 52;
        test_data[347] = 33'd3291818831;
        test_addr[348] = 53;
        test_data[348] = 33'd48823010;
        test_addr[349] = 54;
        test_data[349] = 33'd1614540136;
        test_addr[350] = 55;
        test_data[350] = 33'd4193154773;
        test_addr[351] = 56;
        test_data[351] = 33'd2473651066;
        test_addr[352] = 57;
        test_data[352] = 33'd22011062;
        test_addr[353] = 58;
        test_data[353] = 33'd3203147784;
        test_addr[354] = 59;
        test_data[354] = 33'd1487397129;
        test_addr[355] = 60;
        test_data[355] = 33'd6717228421;
        test_addr[356] = 61;
        test_data[356] = 33'd2535377820;
        test_addr[357] = 62;
        test_data[357] = 33'd504570280;
        test_addr[358] = 63;
        test_data[358] = 33'd7440189888;
        test_addr[359] = 64;
        test_data[359] = 33'd4168218661;
        test_addr[360] = 65;
        test_data[360] = 33'd4169485515;
        test_addr[361] = 160;
        test_data[361] = 33'd2220794859;
        test_addr[362] = 161;
        test_data[362] = 33'd8201736234;
        test_addr[363] = 162;
        test_data[363] = 33'd775522268;
        test_addr[364] = 163;
        test_data[364] = 33'd3495425455;
        test_addr[365] = 164;
        test_data[365] = 33'd2460820341;
        test_addr[366] = 165;
        test_data[366] = 33'd3760476342;
        test_addr[367] = 626;
        test_data[367] = 33'd6482080724;
        test_addr[368] = 627;
        test_data[368] = 33'd2689636519;
        test_addr[369] = 628;
        test_data[369] = 33'd2469942537;
        test_addr[370] = 629;
        test_data[370] = 33'd7627375600;
        test_addr[371] = 630;
        test_data[371] = 33'd3572526873;
        test_addr[372] = 631;
        test_data[372] = 33'd7326789471;
        test_addr[373] = 632;
        test_data[373] = 33'd3201343516;
        test_addr[374] = 633;
        test_data[374] = 33'd1874676766;
        test_addr[375] = 634;
        test_data[375] = 33'd954992338;
        test_addr[376] = 635;
        test_data[376] = 33'd2466428267;
        test_addr[377] = 636;
        test_data[377] = 33'd4218479966;
        test_addr[378] = 637;
        test_data[378] = 33'd8090133021;
        test_addr[379] = 638;
        test_data[379] = 33'd881995127;
        test_addr[380] = 639;
        test_data[380] = 33'd1193599707;
        test_addr[381] = 640;
        test_data[381] = 33'd1559299331;
        test_addr[382] = 641;
        test_data[382] = 33'd2087204287;
        test_addr[383] = 642;
        test_data[383] = 33'd7557932772;
        test_addr[384] = 643;
        test_data[384] = 33'd4156477301;
        test_addr[385] = 644;
        test_data[385] = 33'd3175733827;
        test_addr[386] = 645;
        test_data[386] = 33'd2042867590;
        test_addr[387] = 646;
        test_data[387] = 33'd6032340137;
        test_addr[388] = 647;
        test_data[388] = 33'd3927182985;
        test_addr[389] = 648;
        test_data[389] = 33'd3673972943;
        test_addr[390] = 649;
        test_data[390] = 33'd2151483163;
        test_addr[391] = 650;
        test_data[391] = 33'd8450622538;
        test_addr[392] = 651;
        test_data[392] = 33'd2006915388;
        test_addr[393] = 166;
        test_data[393] = 33'd1889795081;
        test_addr[394] = 167;
        test_data[394] = 33'd3268472177;
        test_addr[395] = 168;
        test_data[395] = 33'd8558962168;
        test_addr[396] = 169;
        test_data[396] = 33'd1140743891;
        test_addr[397] = 170;
        test_data[397] = 33'd3539743854;
        test_addr[398] = 171;
        test_data[398] = 33'd3511614128;
        test_addr[399] = 172;
        test_data[399] = 33'd5954061798;
        test_addr[400] = 173;
        test_data[400] = 33'd422894365;
        test_addr[401] = 174;
        test_data[401] = 33'd7674608762;
        test_addr[402] = 175;
        test_data[402] = 33'd3567745488;
        test_addr[403] = 176;
        test_data[403] = 33'd5381996351;
        test_addr[404] = 177;
        test_data[404] = 33'd2295881178;
        test_addr[405] = 178;
        test_data[405] = 33'd2677761729;
        test_addr[406] = 89;
        test_data[406] = 33'd1036241526;
        test_addr[407] = 90;
        test_data[407] = 33'd548807498;
        test_addr[408] = 91;
        test_data[408] = 33'd3415150818;
        test_addr[409] = 92;
        test_data[409] = 33'd4105109197;
        test_addr[410] = 93;
        test_data[410] = 33'd4579174745;
        test_addr[411] = 94;
        test_data[411] = 33'd2640578934;
        test_addr[412] = 179;
        test_data[412] = 33'd2886227464;
        test_addr[413] = 180;
        test_data[413] = 33'd1980496809;
        test_addr[414] = 181;
        test_data[414] = 33'd3424920418;
        test_addr[415] = 182;
        test_data[415] = 33'd1222529405;
        test_addr[416] = 183;
        test_data[416] = 33'd4192569996;
        test_addr[417] = 184;
        test_data[417] = 33'd961772350;
        test_addr[418] = 185;
        test_data[418] = 33'd8012074517;
        test_addr[419] = 186;
        test_data[419] = 33'd2175561490;
        test_addr[420] = 602;
        test_data[420] = 33'd5519892082;
        test_addr[421] = 603;
        test_data[421] = 33'd434815353;
        test_addr[422] = 604;
        test_data[422] = 33'd152904658;
        test_addr[423] = 605;
        test_data[423] = 33'd4068052147;
        test_addr[424] = 606;
        test_data[424] = 33'd906696308;
        test_addr[425] = 607;
        test_data[425] = 33'd3685335968;
        test_addr[426] = 608;
        test_data[426] = 33'd3635138265;
        test_addr[427] = 609;
        test_data[427] = 33'd7300146947;
        test_addr[428] = 610;
        test_data[428] = 33'd2988230185;
        test_addr[429] = 611;
        test_data[429] = 33'd4475360625;
        test_addr[430] = 612;
        test_data[430] = 33'd2469017315;
        test_addr[431] = 613;
        test_data[431] = 33'd3646976116;
        test_addr[432] = 614;
        test_data[432] = 33'd2005415173;
        test_addr[433] = 615;
        test_data[433] = 33'd5290442024;
        test_addr[434] = 616;
        test_data[434] = 33'd1306428470;
        test_addr[435] = 617;
        test_data[435] = 33'd4082994306;
        test_addr[436] = 618;
        test_data[436] = 33'd902420674;
        test_addr[437] = 619;
        test_data[437] = 33'd8381963636;
        test_addr[438] = 620;
        test_data[438] = 33'd3343656720;
        test_addr[439] = 621;
        test_data[439] = 33'd723470077;
        test_addr[440] = 187;
        test_data[440] = 33'd3131077888;
        test_addr[441] = 188;
        test_data[441] = 33'd128496091;
        test_addr[442] = 189;
        test_data[442] = 33'd133639369;
        test_addr[443] = 190;
        test_data[443] = 33'd4284820396;
        test_addr[444] = 191;
        test_data[444] = 33'd3150765077;
        test_addr[445] = 192;
        test_data[445] = 33'd4570008617;
        test_addr[446] = 193;
        test_data[446] = 33'd4417566192;
        test_addr[447] = 194;
        test_data[447] = 33'd2242595831;
        test_addr[448] = 195;
        test_data[448] = 33'd7536478525;
        test_addr[449] = 196;
        test_data[449] = 33'd1811402878;
        test_addr[450] = 197;
        test_data[450] = 33'd4914750613;
        test_addr[451] = 198;
        test_data[451] = 33'd1771443269;
        test_addr[452] = 199;
        test_data[452] = 33'd1445264864;
        test_addr[453] = 200;
        test_data[453] = 33'd3635105000;
        test_addr[454] = 201;
        test_data[454] = 33'd6217612467;
        test_addr[455] = 202;
        test_data[455] = 33'd4173384693;
        test_addr[456] = 667;
        test_data[456] = 33'd6543946986;
        test_addr[457] = 668;
        test_data[457] = 33'd7105839455;
        test_addr[458] = 669;
        test_data[458] = 33'd879311410;
        test_addr[459] = 670;
        test_data[459] = 33'd7492847092;
        test_addr[460] = 671;
        test_data[460] = 33'd3754236325;
        test_addr[461] = 672;
        test_data[461] = 33'd5706595733;
        test_addr[462] = 673;
        test_data[462] = 33'd1252547980;
        test_addr[463] = 674;
        test_data[463] = 33'd993674477;
        test_addr[464] = 675;
        test_data[464] = 33'd7360008379;
        test_addr[465] = 676;
        test_data[465] = 33'd2458873297;
        test_addr[466] = 677;
        test_data[466] = 33'd3780631796;
        test_addr[467] = 203;
        test_data[467] = 33'd1663091370;
        test_addr[468] = 204;
        test_data[468] = 33'd7929684744;
        test_addr[469] = 205;
        test_data[469] = 33'd349509858;
        test_addr[470] = 206;
        test_data[470] = 33'd871555750;
        test_addr[471] = 207;
        test_data[471] = 33'd3823761644;
        test_addr[472] = 208;
        test_data[472] = 33'd3010632164;
        test_addr[473] = 209;
        test_data[473] = 33'd6396403772;
        test_addr[474] = 210;
        test_data[474] = 33'd2556735740;
        test_addr[475] = 211;
        test_data[475] = 33'd3337632621;
        test_addr[476] = 212;
        test_data[476] = 33'd7272814496;
        test_addr[477] = 213;
        test_data[477] = 33'd371999850;
        test_addr[478] = 214;
        test_data[478] = 33'd3364977113;
        test_addr[479] = 215;
        test_data[479] = 33'd2179149214;
        test_addr[480] = 216;
        test_data[480] = 33'd2231833515;
        test_addr[481] = 217;
        test_data[481] = 33'd797224449;
        test_addr[482] = 218;
        test_data[482] = 33'd2791150383;
        test_addr[483] = 219;
        test_data[483] = 33'd7888938216;
        test_addr[484] = 220;
        test_data[484] = 33'd4233481341;
        test_addr[485] = 221;
        test_data[485] = 33'd285286831;
        test_addr[486] = 222;
        test_data[486] = 33'd8528701038;
        test_addr[487] = 222;
        test_data[487] = 33'd4233733742;
        test_addr[488] = 223;
        test_data[488] = 33'd308136402;
        test_addr[489] = 224;
        test_data[489] = 33'd6438596732;
        test_addr[490] = 223;
        test_data[490] = 33'd308136402;
        test_addr[491] = 224;
        test_data[491] = 33'd2143629436;
        test_addr[492] = 225;
        test_data[492] = 33'd5550779402;
        test_addr[493] = 226;
        test_data[493] = 33'd5687314748;
        test_addr[494] = 227;
        test_data[494] = 33'd5314626400;
        test_addr[495] = 228;
        test_data[495] = 33'd7113987233;
        test_addr[496] = 830;
        test_data[496] = 33'd72105947;
        test_addr[497] = 831;
        test_data[497] = 33'd8261219150;
        test_addr[498] = 832;
        test_data[498] = 33'd4001181699;
        test_addr[499] = 833;
        test_data[499] = 33'd1217572098;
        test_addr[500] = 834;
        test_data[500] = 33'd4233557749;
        test_addr[501] = 835;
        test_data[501] = 33'd4756690905;
        test_addr[502] = 836;
        test_data[502] = 33'd4728319758;
        test_addr[503] = 229;
        test_data[503] = 33'd5140199940;
        test_addr[504] = 230;
        test_data[504] = 33'd4387034904;
        test_addr[505] = 231;
        test_data[505] = 33'd1221449456;
        test_addr[506] = 946;
        test_data[506] = 33'd1984305920;
        test_addr[507] = 947;
        test_data[507] = 33'd7692639235;
        test_addr[508] = 948;
        test_data[508] = 33'd4984941441;
        test_addr[509] = 232;
        test_data[509] = 33'd4110523392;
        test_addr[510] = 233;
        test_data[510] = 33'd2577766004;
        test_addr[511] = 234;
        test_data[511] = 33'd5040390600;
        test_addr[512] = 937;
        test_data[512] = 33'd625389764;
        test_addr[513] = 938;
        test_data[513] = 33'd8217814515;
        test_addr[514] = 939;
        test_data[514] = 33'd8557709683;
        test_addr[515] = 940;
        test_data[515] = 33'd3211187226;
        test_addr[516] = 941;
        test_data[516] = 33'd1873325343;
        test_addr[517] = 942;
        test_data[517] = 33'd3185997769;
        test_addr[518] = 943;
        test_data[518] = 33'd1653503808;
        test_addr[519] = 944;
        test_data[519] = 33'd1934668787;
        test_addr[520] = 945;
        test_data[520] = 33'd1578395060;
        test_addr[521] = 946;
        test_data[521] = 33'd1984305920;
        test_addr[522] = 947;
        test_data[522] = 33'd3397671939;
        test_addr[523] = 948;
        test_data[523] = 33'd689974145;
        test_addr[524] = 949;
        test_data[524] = 33'd1182899197;
        test_addr[525] = 950;
        test_data[525] = 33'd2459752245;
        test_addr[526] = 951;
        test_data[526] = 33'd3631193825;
        test_addr[527] = 952;
        test_data[527] = 33'd1791314849;
        test_addr[528] = 953;
        test_data[528] = 33'd2693867941;
        test_addr[529] = 954;
        test_data[529] = 33'd7091615423;
        test_addr[530] = 955;
        test_data[530] = 33'd905894982;
        test_addr[531] = 956;
        test_data[531] = 33'd90020364;
        test_addr[532] = 957;
        test_data[532] = 33'd2991872276;
        test_addr[533] = 958;
        test_data[533] = 33'd3447221745;
        test_addr[534] = 959;
        test_data[534] = 33'd1132988677;
        test_addr[535] = 960;
        test_data[535] = 33'd7792132987;
        test_addr[536] = 961;
        test_data[536] = 33'd6370015393;
        test_addr[537] = 962;
        test_data[537] = 33'd2765447673;
        test_addr[538] = 963;
        test_data[538] = 33'd6451783245;
        test_addr[539] = 964;
        test_data[539] = 33'd3129425578;
        test_addr[540] = 965;
        test_data[540] = 33'd6679131125;
        test_addr[541] = 966;
        test_data[541] = 33'd2560894838;
        test_addr[542] = 967;
        test_data[542] = 33'd2075372781;
        test_addr[543] = 968;
        test_data[543] = 33'd7369061236;
        test_addr[544] = 969;
        test_data[544] = 33'd6248436800;
        test_addr[545] = 970;
        test_data[545] = 33'd4208904194;
        test_addr[546] = 971;
        test_data[546] = 33'd1365898262;
        test_addr[547] = 972;
        test_data[547] = 33'd1158453115;
        test_addr[548] = 973;
        test_data[548] = 33'd3512163126;
        test_addr[549] = 974;
        test_data[549] = 33'd1819208149;
        test_addr[550] = 975;
        test_data[550] = 33'd900993035;
        test_addr[551] = 976;
        test_data[551] = 33'd888555328;
        test_addr[552] = 977;
        test_data[552] = 33'd871000283;
        test_addr[553] = 978;
        test_data[553] = 33'd1143928461;
        test_addr[554] = 979;
        test_data[554] = 33'd3552257411;
        test_addr[555] = 980;
        test_data[555] = 33'd8016854113;
        test_addr[556] = 981;
        test_data[556] = 33'd4301773313;
        test_addr[557] = 982;
        test_data[557] = 33'd6359390204;
        test_addr[558] = 235;
        test_data[558] = 33'd1995153683;
        test_addr[559] = 494;
        test_data[559] = 33'd6841726114;
        test_addr[560] = 495;
        test_data[560] = 33'd1266991624;
        test_addr[561] = 496;
        test_data[561] = 33'd1858394599;
        test_addr[562] = 497;
        test_data[562] = 33'd2724175409;
        test_addr[563] = 498;
        test_data[563] = 33'd5614661622;
        test_addr[564] = 236;
        test_data[564] = 33'd3308823479;
        test_addr[565] = 237;
        test_data[565] = 33'd3710833553;
        test_addr[566] = 238;
        test_data[566] = 33'd5833139424;
        test_addr[567] = 239;
        test_data[567] = 33'd5275264421;
        test_addr[568] = 240;
        test_data[568] = 33'd2785262700;
        test_addr[569] = 241;
        test_data[569] = 33'd3647911902;
        test_addr[570] = 242;
        test_data[570] = 33'd1066521417;
        test_addr[571] = 243;
        test_data[571] = 33'd488961057;
        test_addr[572] = 244;
        test_data[572] = 33'd2896346636;
        test_addr[573] = 245;
        test_data[573] = 33'd2801824671;
        test_addr[574] = 246;
        test_data[574] = 33'd2321687399;
        test_addr[575] = 247;
        test_data[575] = 33'd2088915050;
        test_addr[576] = 248;
        test_data[576] = 33'd2567675747;
        test_addr[577] = 249;
        test_data[577] = 33'd634363534;
        test_addr[578] = 250;
        test_data[578] = 33'd3563604010;
        test_addr[579] = 251;
        test_data[579] = 33'd528276894;
        test_addr[580] = 969;
        test_data[580] = 33'd1953469504;
        test_addr[581] = 252;
        test_data[581] = 33'd3233104755;
        test_addr[582] = 253;
        test_data[582] = 33'd2251486923;
        test_addr[583] = 254;
        test_data[583] = 33'd4129721780;
        test_addr[584] = 255;
        test_data[584] = 33'd5908754263;
        test_addr[585] = 256;
        test_data[585] = 33'd214161842;
        test_addr[586] = 257;
        test_data[586] = 33'd7055571207;
        test_addr[587] = 258;
        test_data[587] = 33'd3768261454;
        test_addr[588] = 259;
        test_data[588] = 33'd735052196;
        test_addr[589] = 260;
        test_data[589] = 33'd2209658087;
        test_addr[590] = 261;
        test_data[590] = 33'd2908678289;
        test_addr[591] = 262;
        test_data[591] = 33'd3668048787;
        test_addr[592] = 263;
        test_data[592] = 33'd2095898228;
        test_addr[593] = 264;
        test_data[593] = 33'd1563802891;
        test_addr[594] = 265;
        test_data[594] = 33'd6493953492;
        test_addr[595] = 266;
        test_data[595] = 33'd247106196;
        test_addr[596] = 267;
        test_data[596] = 33'd1193893598;
        test_addr[597] = 268;
        test_data[597] = 33'd458908171;
        test_addr[598] = 269;
        test_data[598] = 33'd7589653210;
        test_addr[599] = 270;
        test_data[599] = 33'd1805982290;
        test_addr[600] = 271;
        test_data[600] = 33'd2912190139;
        test_addr[601] = 272;
        test_data[601] = 33'd495494873;
        test_addr[602] = 273;
        test_data[602] = 33'd5558780609;
        test_addr[603] = 274;
        test_data[603] = 33'd5769817226;
        test_addr[604] = 92;
        test_data[604] = 33'd4105109197;
        test_addr[605] = 93;
        test_data[605] = 33'd284207449;
        test_addr[606] = 94;
        test_data[606] = 33'd2640578934;
        test_addr[607] = 95;
        test_data[607] = 33'd5062083936;
        test_addr[608] = 96;
        test_data[608] = 33'd5735974740;
        test_addr[609] = 97;
        test_data[609] = 33'd2681259618;
        test_addr[610] = 98;
        test_data[610] = 33'd1885671812;
        test_addr[611] = 99;
        test_data[611] = 33'd2668054470;
        test_addr[612] = 100;
        test_data[612] = 33'd7368675152;
        test_addr[613] = 101;
        test_data[613] = 33'd1530703461;
        test_addr[614] = 275;
        test_data[614] = 33'd94646178;
        test_addr[615] = 276;
        test_data[615] = 33'd3369498205;
        test_addr[616] = 277;
        test_data[616] = 33'd76492403;
        test_addr[617] = 278;
        test_data[617] = 33'd7779739427;
        test_addr[618] = 279;
        test_data[618] = 33'd1301179723;
        test_addr[619] = 280;
        test_data[619] = 33'd535207050;
        test_addr[620] = 281;
        test_data[620] = 33'd7400389074;
        test_addr[621] = 282;
        test_data[621] = 33'd1396158732;
        test_addr[622] = 283;
        test_data[622] = 33'd4134955926;
        test_addr[623] = 284;
        test_data[623] = 33'd1470833253;
        test_addr[624] = 417;
        test_data[624] = 33'd3832011826;
        test_addr[625] = 418;
        test_data[625] = 33'd1591263160;
        test_addr[626] = 419;
        test_data[626] = 33'd188335908;
        test_addr[627] = 420;
        test_data[627] = 33'd4738805490;
        test_addr[628] = 421;
        test_data[628] = 33'd3567358548;
        test_addr[629] = 422;
        test_data[629] = 33'd2973342047;
        test_addr[630] = 423;
        test_data[630] = 33'd5968912572;
        test_addr[631] = 424;
        test_data[631] = 33'd458707520;
        test_addr[632] = 425;
        test_data[632] = 33'd6639308970;
        test_addr[633] = 426;
        test_data[633] = 33'd138557177;
        test_addr[634] = 427;
        test_data[634] = 33'd1979928705;
        test_addr[635] = 428;
        test_data[635] = 33'd1479974522;
        test_addr[636] = 429;
        test_data[636] = 33'd3385333427;
        test_addr[637] = 430;
        test_data[637] = 33'd2489047385;
        test_addr[638] = 431;
        test_data[638] = 33'd723449661;
        test_addr[639] = 432;
        test_data[639] = 33'd1474827311;
        test_addr[640] = 433;
        test_data[640] = 33'd5039391830;
        test_addr[641] = 434;
        test_data[641] = 33'd3881600915;
        test_addr[642] = 435;
        test_data[642] = 33'd1781223650;
        test_addr[643] = 436;
        test_data[643] = 33'd1024435444;
        test_addr[644] = 437;
        test_data[644] = 33'd4685483373;
        test_addr[645] = 438;
        test_data[645] = 33'd3957892093;
        test_addr[646] = 439;
        test_data[646] = 33'd4682735552;
        test_addr[647] = 440;
        test_data[647] = 33'd118271122;
        test_addr[648] = 285;
        test_data[648] = 33'd7984929193;
        test_addr[649] = 286;
        test_data[649] = 33'd1109364526;
        test_addr[650] = 287;
        test_data[650] = 33'd2077233220;
        test_addr[651] = 288;
        test_data[651] = 33'd3761039539;
        test_addr[652] = 289;
        test_data[652] = 33'd940573815;
        test_addr[653] = 290;
        test_data[653] = 33'd1919999915;
        test_addr[654] = 291;
        test_data[654] = 33'd2648754452;
        test_addr[655] = 292;
        test_data[655] = 33'd3646512956;
        test_addr[656] = 293;
        test_data[656] = 33'd120765790;
        test_addr[657] = 294;
        test_data[657] = 33'd6652519248;
        test_addr[658] = 295;
        test_data[658] = 33'd431105951;
        test_addr[659] = 296;
        test_data[659] = 33'd8208403991;
        test_addr[660] = 297;
        test_data[660] = 33'd7488600754;
        test_addr[661] = 141;
        test_data[661] = 33'd3385276041;
        test_addr[662] = 142;
        test_data[662] = 33'd2889759130;
        test_addr[663] = 143;
        test_data[663] = 33'd6218250061;
        test_addr[664] = 144;
        test_data[664] = 33'd3584443635;
        test_addr[665] = 145;
        test_data[665] = 33'd2276121759;
        test_addr[666] = 146;
        test_data[666] = 33'd1978812597;
        test_addr[667] = 147;
        test_data[667] = 33'd3498313420;
        test_addr[668] = 148;
        test_data[668] = 33'd4014633640;
        test_addr[669] = 149;
        test_data[669] = 33'd4309978280;
        test_addr[670] = 150;
        test_data[670] = 33'd1729930243;
        test_addr[671] = 151;
        test_data[671] = 33'd4477946697;
        test_addr[672] = 152;
        test_data[672] = 33'd7654255503;
        test_addr[673] = 153;
        test_data[673] = 33'd352254805;
        test_addr[674] = 154;
        test_data[674] = 33'd6682840204;
        test_addr[675] = 155;
        test_data[675] = 33'd979919250;
        test_addr[676] = 156;
        test_data[676] = 33'd1324821377;
        test_addr[677] = 157;
        test_data[677] = 33'd6385333335;
        test_addr[678] = 158;
        test_data[678] = 33'd2395849516;
        test_addr[679] = 298;
        test_data[679] = 33'd3316398040;
        test_addr[680] = 299;
        test_data[680] = 33'd1285349339;
        test_addr[681] = 300;
        test_data[681] = 33'd4260493041;
        test_addr[682] = 301;
        test_data[682] = 33'd779647779;
        test_addr[683] = 302;
        test_data[683] = 33'd2759854552;
        test_addr[684] = 303;
        test_data[684] = 33'd4718411272;
        test_addr[685] = 304;
        test_data[685] = 33'd6300220529;
        test_addr[686] = 305;
        test_data[686] = 33'd6161202446;
        test_addr[687] = 306;
        test_data[687] = 33'd1400119106;
        test_addr[688] = 713;
        test_data[688] = 33'd3261845956;
        test_addr[689] = 714;
        test_data[689] = 33'd4226705526;
        test_addr[690] = 715;
        test_data[690] = 33'd3264214500;
        test_addr[691] = 716;
        test_data[691] = 33'd3183387761;
        test_addr[692] = 717;
        test_data[692] = 33'd3532130073;
        test_addr[693] = 718;
        test_data[693] = 33'd2494614555;
        test_addr[694] = 719;
        test_data[694] = 33'd6743677968;
        test_addr[695] = 720;
        test_data[695] = 33'd2104937406;
        test_addr[696] = 721;
        test_data[696] = 33'd2025627376;
        test_addr[697] = 722;
        test_data[697] = 33'd6952921341;
        test_addr[698] = 723;
        test_data[698] = 33'd3748128516;
        test_addr[699] = 724;
        test_data[699] = 33'd7859574700;
        test_addr[700] = 725;
        test_data[700] = 33'd3136553366;
        test_addr[701] = 726;
        test_data[701] = 33'd1207862729;
        test_addr[702] = 307;
        test_data[702] = 33'd3130498011;
        test_addr[703] = 282;
        test_data[703] = 33'd1396158732;
        test_addr[704] = 283;
        test_data[704] = 33'd4134955926;
        test_addr[705] = 284;
        test_data[705] = 33'd1470833253;
        test_addr[706] = 285;
        test_data[706] = 33'd3689961897;
        test_addr[707] = 286;
        test_data[707] = 33'd1109364526;
        test_addr[708] = 287;
        test_data[708] = 33'd2077233220;
        test_addr[709] = 288;
        test_data[709] = 33'd8322104245;
        test_addr[710] = 289;
        test_data[710] = 33'd940573815;
        test_addr[711] = 290;
        test_data[711] = 33'd7240485132;
        test_addr[712] = 308;
        test_data[712] = 33'd2611705428;
        test_addr[713] = 309;
        test_data[713] = 33'd3941608837;
        test_addr[714] = 310;
        test_data[714] = 33'd3094631771;
        test_addr[715] = 311;
        test_data[715] = 33'd1449524691;
        test_addr[716] = 312;
        test_data[716] = 33'd240548675;
        test_addr[717] = 313;
        test_data[717] = 33'd3069166694;
        test_addr[718] = 314;
        test_data[718] = 33'd6436033102;
        test_addr[719] = 315;
        test_data[719] = 33'd3309303920;
        test_addr[720] = 316;
        test_data[720] = 33'd7053424836;
        test_addr[721] = 317;
        test_data[721] = 33'd4112356272;
        test_addr[722] = 318;
        test_data[722] = 33'd1367187386;
        test_addr[723] = 319;
        test_data[723] = 33'd398366425;
        test_addr[724] = 320;
        test_data[724] = 33'd2213105581;
        test_addr[725] = 321;
        test_data[725] = 33'd4078285937;
        test_addr[726] = 724;
        test_data[726] = 33'd3564607404;
        test_addr[727] = 725;
        test_data[727] = 33'd3136553366;
        test_addr[728] = 726;
        test_data[728] = 33'd1207862729;
        test_addr[729] = 727;
        test_data[729] = 33'd1005793312;
        test_addr[730] = 728;
        test_data[730] = 33'd5579284531;
        test_addr[731] = 729;
        test_data[731] = 33'd5214312842;
        test_addr[732] = 730;
        test_data[732] = 33'd8362896084;
        test_addr[733] = 731;
        test_data[733] = 33'd1353510671;
        test_addr[734] = 732;
        test_data[734] = 33'd7833717569;
        test_addr[735] = 733;
        test_data[735] = 33'd1312293725;
        test_addr[736] = 734;
        test_data[736] = 33'd7447473199;
        test_addr[737] = 735;
        test_data[737] = 33'd567958459;
        test_addr[738] = 736;
        test_data[738] = 33'd5219266647;
        test_addr[739] = 737;
        test_data[739] = 33'd7665912340;
        test_addr[740] = 738;
        test_data[740] = 33'd791004845;
        test_addr[741] = 739;
        test_data[741] = 33'd3426545964;
        test_addr[742] = 740;
        test_data[742] = 33'd7528115033;
        test_addr[743] = 741;
        test_data[743] = 33'd1810153704;
        test_addr[744] = 742;
        test_data[744] = 33'd2878401245;
        test_addr[745] = 743;
        test_data[745] = 33'd6785677295;
        test_addr[746] = 744;
        test_data[746] = 33'd7509780377;
        test_addr[747] = 745;
        test_data[747] = 33'd3435630877;
        test_addr[748] = 746;
        test_data[748] = 33'd3185922216;
        test_addr[749] = 747;
        test_data[749] = 33'd7696572917;
        test_addr[750] = 748;
        test_data[750] = 33'd5816797086;
        test_addr[751] = 749;
        test_data[751] = 33'd1248251572;
        test_addr[752] = 750;
        test_data[752] = 33'd282558174;
        test_addr[753] = 751;
        test_data[753] = 33'd3419461017;
        test_addr[754] = 752;
        test_data[754] = 33'd467983000;
        test_addr[755] = 753;
        test_data[755] = 33'd8396447271;
        test_addr[756] = 754;
        test_data[756] = 33'd2930249500;
        test_addr[757] = 755;
        test_data[757] = 33'd4522075247;
        test_addr[758] = 756;
        test_data[758] = 33'd5632998267;
        test_addr[759] = 322;
        test_data[759] = 33'd4172724571;
        test_addr[760] = 323;
        test_data[760] = 33'd2407757486;
        test_addr[761] = 324;
        test_data[761] = 33'd2439471225;
        test_addr[762] = 325;
        test_data[762] = 33'd2995637218;
        test_addr[763] = 326;
        test_data[763] = 33'd4825498686;
        test_addr[764] = 327;
        test_data[764] = 33'd318989378;
        test_addr[765] = 328;
        test_data[765] = 33'd3131202390;
        test_addr[766] = 329;
        test_data[766] = 33'd7434815525;
        test_addr[767] = 330;
        test_data[767] = 33'd1703867803;
        test_addr[768] = 331;
        test_data[768] = 33'd2887064224;
        test_addr[769] = 332;
        test_data[769] = 33'd6677737118;
        test_addr[770] = 333;
        test_data[770] = 33'd1462324255;
        test_addr[771] = 334;
        test_data[771] = 33'd3909284796;
        test_addr[772] = 335;
        test_data[772] = 33'd115410482;
        test_addr[773] = 336;
        test_data[773] = 33'd2188727585;
        test_addr[774] = 337;
        test_data[774] = 33'd6461955697;
        test_addr[775] = 338;
        test_data[775] = 33'd3556465203;
        test_addr[776] = 865;
        test_data[776] = 33'd3049915918;
        test_addr[777] = 866;
        test_data[777] = 33'd2528451676;
        test_addr[778] = 867;
        test_data[778] = 33'd4195620311;
        test_addr[779] = 339;
        test_data[779] = 33'd6682629276;
        test_addr[780] = 340;
        test_data[780] = 33'd4746381244;
        test_addr[781] = 341;
        test_data[781] = 33'd829190514;
        test_addr[782] = 342;
        test_data[782] = 33'd2723057950;
        test_addr[783] = 343;
        test_data[783] = 33'd1636516063;
        test_addr[784] = 39;
        test_data[784] = 33'd4629947426;
        test_addr[785] = 40;
        test_data[785] = 33'd5005863210;
        test_addr[786] = 41;
        test_data[786] = 33'd6799980467;
        test_addr[787] = 42;
        test_data[787] = 33'd8409078549;
        test_addr[788] = 43;
        test_data[788] = 33'd1598694208;
        test_addr[789] = 44;
        test_data[789] = 33'd498645939;
        test_addr[790] = 45;
        test_data[790] = 33'd2757741745;
        test_addr[791] = 46;
        test_data[791] = 33'd317333202;
        test_addr[792] = 47;
        test_data[792] = 33'd4813649833;
        test_addr[793] = 48;
        test_data[793] = 33'd2577690104;
        test_addr[794] = 344;
        test_data[794] = 33'd281373290;
        test_addr[795] = 251;
        test_data[795] = 33'd4941625912;
        test_addr[796] = 252;
        test_data[796] = 33'd3233104755;
        test_addr[797] = 253;
        test_data[797] = 33'd2251486923;
        test_addr[798] = 254;
        test_data[798] = 33'd4129721780;
        test_addr[799] = 255;
        test_data[799] = 33'd1613786967;
        test_addr[800] = 256;
        test_data[800] = 33'd214161842;
        test_addr[801] = 257;
        test_data[801] = 33'd2760603911;
        test_addr[802] = 258;
        test_data[802] = 33'd3768261454;
        test_addr[803] = 259;
        test_data[803] = 33'd5698584015;
        test_addr[804] = 260;
        test_data[804] = 33'd2209658087;
        test_addr[805] = 261;
        test_data[805] = 33'd2908678289;
        test_addr[806] = 262;
        test_data[806] = 33'd3668048787;
        test_addr[807] = 263;
        test_data[807] = 33'd2095898228;
        test_addr[808] = 264;
        test_data[808] = 33'd1563802891;
        test_addr[809] = 265;
        test_data[809] = 33'd2198986196;
        test_addr[810] = 266;
        test_data[810] = 33'd247106196;
        test_addr[811] = 267;
        test_data[811] = 33'd8115508662;
        test_addr[812] = 268;
        test_data[812] = 33'd458908171;
        test_addr[813] = 269;
        test_data[813] = 33'd4418602691;
        test_addr[814] = 270;
        test_data[814] = 33'd1805982290;
        test_addr[815] = 271;
        test_data[815] = 33'd6730967967;
        test_addr[816] = 345;
        test_data[816] = 33'd3249490296;
        test_addr[817] = 346;
        test_data[817] = 33'd4865991968;
        test_addr[818] = 347;
        test_data[818] = 33'd184952467;
        test_addr[819] = 348;
        test_data[819] = 33'd7927001949;
        test_addr[820] = 349;
        test_data[820] = 33'd516820221;
        test_addr[821] = 350;
        test_data[821] = 33'd1118902313;
        test_addr[822] = 351;
        test_data[822] = 33'd5372619417;
        test_addr[823] = 352;
        test_data[823] = 33'd147931898;
        test_addr[824] = 353;
        test_data[824] = 33'd5844231282;
        test_addr[825] = 354;
        test_data[825] = 33'd3966319412;
        test_addr[826] = 355;
        test_data[826] = 33'd3274769757;
        test_addr[827] = 356;
        test_data[827] = 33'd5658381331;
        test_addr[828] = 357;
        test_data[828] = 33'd8431968778;
        test_addr[829] = 358;
        test_data[829] = 33'd928067253;
        test_addr[830] = 359;
        test_data[830] = 33'd4082684122;
        test_addr[831] = 360;
        test_data[831] = 33'd5972009549;
        test_addr[832] = 361;
        test_data[832] = 33'd851421913;
        test_addr[833] = 362;
        test_data[833] = 33'd5034836920;
        test_addr[834] = 363;
        test_data[834] = 33'd7739254264;
        test_addr[835] = 364;
        test_data[835] = 33'd4047546126;
        test_addr[836] = 365;
        test_data[836] = 33'd5303177410;
        test_addr[837] = 366;
        test_data[837] = 33'd2115114658;
        test_addr[838] = 367;
        test_data[838] = 33'd916394114;
        test_addr[839] = 368;
        test_data[839] = 33'd5845836600;
        test_addr[840] = 369;
        test_data[840] = 33'd6475150932;
        test_addr[841] = 370;
        test_data[841] = 33'd2827239166;
        test_addr[842] = 588;
        test_data[842] = 33'd1893529001;
        test_addr[843] = 589;
        test_data[843] = 33'd7809953208;
        test_addr[844] = 590;
        test_data[844] = 33'd2083229337;
        test_addr[845] = 591;
        test_data[845] = 33'd4756732875;
        test_addr[846] = 371;
        test_data[846] = 33'd6091737777;
        test_addr[847] = 372;
        test_data[847] = 33'd3348876813;
        test_addr[848] = 373;
        test_data[848] = 33'd6943526;
        test_addr[849] = 374;
        test_data[849] = 33'd6132151847;
        test_addr[850] = 165;
        test_data[850] = 33'd3760476342;
        test_addr[851] = 166;
        test_data[851] = 33'd1889795081;
        test_addr[852] = 167;
        test_data[852] = 33'd6231215534;
        test_addr[853] = 168;
        test_data[853] = 33'd4263994872;
        test_addr[854] = 169;
        test_data[854] = 33'd1140743891;
        test_addr[855] = 375;
        test_data[855] = 33'd137070870;
        test_addr[856] = 376;
        test_data[856] = 33'd3383574487;
        test_addr[857] = 377;
        test_data[857] = 33'd258678087;
        test_addr[858] = 378;
        test_data[858] = 33'd1707274193;
        test_addr[859] = 932;
        test_data[859] = 33'd572260113;
        test_addr[860] = 933;
        test_data[860] = 33'd4465076143;
        test_addr[861] = 934;
        test_data[861] = 33'd5398174937;
        test_addr[862] = 935;
        test_data[862] = 33'd2013495484;
        test_addr[863] = 936;
        test_data[863] = 33'd607348316;
        test_addr[864] = 937;
        test_data[864] = 33'd625389764;
        test_addr[865] = 938;
        test_data[865] = 33'd3922847219;
        test_addr[866] = 939;
        test_data[866] = 33'd4644599356;
        test_addr[867] = 940;
        test_data[867] = 33'd3211187226;
        test_addr[868] = 941;
        test_data[868] = 33'd5755655908;
        test_addr[869] = 942;
        test_data[869] = 33'd3185997769;
        test_addr[870] = 943;
        test_data[870] = 33'd1653503808;
        test_addr[871] = 944;
        test_data[871] = 33'd1934668787;
        test_addr[872] = 945;
        test_data[872] = 33'd1578395060;
        test_addr[873] = 379;
        test_data[873] = 33'd76696075;
        test_addr[874] = 380;
        test_data[874] = 33'd4157069748;
        test_addr[875] = 381;
        test_data[875] = 33'd3760007301;
        test_addr[876] = 382;
        test_data[876] = 33'd8022734404;
        test_addr[877] = 383;
        test_data[877] = 33'd6328845626;
        test_addr[878] = 384;
        test_data[878] = 33'd7737688341;
        test_addr[879] = 385;
        test_data[879] = 33'd2580136147;
        test_addr[880] = 251;
        test_data[880] = 33'd646658616;
        test_addr[881] = 252;
        test_data[881] = 33'd3233104755;
        test_addr[882] = 253;
        test_data[882] = 33'd2251486923;
        test_addr[883] = 254;
        test_data[883] = 33'd4376600487;
        test_addr[884] = 255;
        test_data[884] = 33'd1613786967;
        test_addr[885] = 256;
        test_data[885] = 33'd214161842;
        test_addr[886] = 257;
        test_data[886] = 33'd6410338394;
        test_addr[887] = 258;
        test_data[887] = 33'd3768261454;
        test_addr[888] = 259;
        test_data[888] = 33'd1403616719;
        test_addr[889] = 260;
        test_data[889] = 33'd2209658087;
        test_addr[890] = 261;
        test_data[890] = 33'd2908678289;
        test_addr[891] = 262;
        test_data[891] = 33'd3668048787;
        test_addr[892] = 263;
        test_data[892] = 33'd2095898228;
        test_addr[893] = 264;
        test_data[893] = 33'd1563802891;
        test_addr[894] = 265;
        test_data[894] = 33'd2198986196;
        test_addr[895] = 266;
        test_data[895] = 33'd247106196;
        test_addr[896] = 267;
        test_data[896] = 33'd3820541366;
        test_addr[897] = 268;
        test_data[897] = 33'd458908171;
        test_addr[898] = 269;
        test_data[898] = 33'd123635395;
        test_addr[899] = 270;
        test_data[899] = 33'd6998582653;
        test_addr[900] = 271;
        test_data[900] = 33'd8302108293;
        test_addr[901] = 272;
        test_data[901] = 33'd495494873;
        test_addr[902] = 386;
        test_data[902] = 33'd2578070289;
        test_addr[903] = 387;
        test_data[903] = 33'd7447882809;
        test_addr[904] = 388;
        test_data[904] = 33'd2217298716;
        test_addr[905] = 389;
        test_data[905] = 33'd2233888802;
        test_addr[906] = 390;
        test_data[906] = 33'd8242931389;
        test_addr[907] = 391;
        test_data[907] = 33'd4156755592;
        test_addr[908] = 392;
        test_data[908] = 33'd4188547242;
        test_addr[909] = 393;
        test_data[909] = 33'd7879783511;
        test_addr[910] = 394;
        test_data[910] = 33'd7815638482;
        test_addr[911] = 448;
        test_data[911] = 33'd4199406484;
        test_addr[912] = 449;
        test_data[912] = 33'd2000661367;
        test_addr[913] = 450;
        test_data[913] = 33'd1220832376;
        test_addr[914] = 451;
        test_data[914] = 33'd2278524113;
        test_addr[915] = 452;
        test_data[915] = 33'd8231868362;
        test_addr[916] = 453;
        test_data[916] = 33'd6910392892;
        test_addr[917] = 454;
        test_data[917] = 33'd6912630279;
        test_addr[918] = 455;
        test_data[918] = 33'd3799628466;
        test_addr[919] = 456;
        test_data[919] = 33'd1297742875;
        test_addr[920] = 457;
        test_data[920] = 33'd2700525639;
        test_addr[921] = 458;
        test_data[921] = 33'd1845881788;
        test_addr[922] = 459;
        test_data[922] = 33'd582707416;
        test_addr[923] = 460;
        test_data[923] = 33'd3277373807;
        test_addr[924] = 395;
        test_data[924] = 33'd6584197819;
        test_addr[925] = 396;
        test_data[925] = 33'd179786261;
        test_addr[926] = 397;
        test_data[926] = 33'd7913683884;
        test_addr[927] = 398;
        test_data[927] = 33'd6419553419;
        test_addr[928] = 399;
        test_data[928] = 33'd3647612275;
        test_addr[929] = 400;
        test_data[929] = 33'd7082142654;
        test_addr[930] = 401;
        test_data[930] = 33'd4710740644;
        test_addr[931] = 402;
        test_data[931] = 33'd246986956;
        test_addr[932] = 403;
        test_data[932] = 33'd4898865076;
        test_addr[933] = 404;
        test_data[933] = 33'd284306586;
        test_addr[934] = 405;
        test_data[934] = 33'd411101395;
        test_addr[935] = 406;
        test_data[935] = 33'd2569288348;
        test_addr[936] = 401;
        test_data[936] = 33'd415773348;
        test_addr[937] = 402;
        test_data[937] = 33'd246986956;
        test_addr[938] = 403;
        test_data[938] = 33'd603897780;
        test_addr[939] = 404;
        test_data[939] = 33'd284306586;
        test_addr[940] = 405;
        test_data[940] = 33'd411101395;
        test_addr[941] = 406;
        test_data[941] = 33'd7125608935;
        test_addr[942] = 407;
        test_data[942] = 33'd4569563985;
        test_addr[943] = 408;
        test_data[943] = 33'd543094332;
        test_addr[944] = 409;
        test_data[944] = 33'd2882373882;
        test_addr[945] = 410;
        test_data[945] = 33'd3422075366;
        test_addr[946] = 411;
        test_data[946] = 33'd7921094178;
        test_addr[947] = 412;
        test_data[947] = 33'd35661170;
        test_addr[948] = 413;
        test_data[948] = 33'd6777784285;
        test_addr[949] = 407;
        test_data[949] = 33'd6802632452;
        test_addr[950] = 408;
        test_data[950] = 33'd543094332;
        test_addr[951] = 409;
        test_data[951] = 33'd2882373882;
        test_addr[952] = 410;
        test_data[952] = 33'd3422075366;
        test_addr[953] = 411;
        test_data[953] = 33'd3626126882;
        test_addr[954] = 412;
        test_data[954] = 33'd35661170;
        test_addr[955] = 169;
        test_data[955] = 33'd6947588909;
        test_addr[956] = 170;
        test_data[956] = 33'd7144715069;
        test_addr[957] = 171;
        test_data[957] = 33'd3511614128;
        test_addr[958] = 172;
        test_data[958] = 33'd1659094502;
        test_addr[959] = 173;
        test_data[959] = 33'd422894365;
        test_addr[960] = 174;
        test_data[960] = 33'd5520444580;
        test_addr[961] = 175;
        test_data[961] = 33'd3567745488;
        test_addr[962] = 176;
        test_data[962] = 33'd1087029055;
        test_addr[963] = 177;
        test_data[963] = 33'd2295881178;
        test_addr[964] = 178;
        test_data[964] = 33'd2677761729;
        test_addr[965] = 179;
        test_data[965] = 33'd2886227464;
        test_addr[966] = 180;
        test_data[966] = 33'd8535352136;
        test_addr[967] = 181;
        test_data[967] = 33'd6492762732;
        test_addr[968] = 182;
        test_data[968] = 33'd1222529405;
        test_addr[969] = 413;
        test_data[969] = 33'd2482816989;
        test_addr[970] = 414;
        test_data[970] = 33'd3438809741;
        test_addr[971] = 415;
        test_data[971] = 33'd2824809495;
        test_addr[972] = 416;
        test_data[972] = 33'd7113925170;
        test_addr[973] = 417;
        test_data[973] = 33'd3832011826;
        test_addr[974] = 61;
        test_data[974] = 33'd6504063154;
        test_addr[975] = 62;
        test_data[975] = 33'd504570280;
        test_addr[976] = 63;
        test_data[976] = 33'd3145222592;
        test_addr[977] = 64;
        test_data[977] = 33'd4168218661;
        test_addr[978] = 65;
        test_data[978] = 33'd4169485515;
        test_addr[979] = 66;
        test_data[979] = 33'd8090029040;
        test_addr[980] = 67;
        test_data[980] = 33'd7076966849;
        test_addr[981] = 68;
        test_data[981] = 33'd2440392340;
        test_addr[982] = 69;
        test_data[982] = 33'd712353462;
        test_addr[983] = 70;
        test_data[983] = 33'd3874690545;
        test_addr[984] = 71;
        test_data[984] = 33'd1800624896;
        test_addr[985] = 72;
        test_data[985] = 33'd3745474962;
        test_addr[986] = 73;
        test_data[986] = 33'd8140864486;
        test_addr[987] = 74;
        test_data[987] = 33'd5490828904;
        test_addr[988] = 75;
        test_data[988] = 33'd3972422453;
        test_addr[989] = 76;
        test_data[989] = 33'd1051232611;
        test_addr[990] = 77;
        test_data[990] = 33'd998193764;
        test_addr[991] = 78;
        test_data[991] = 33'd3591490314;
        test_addr[992] = 79;
        test_data[992] = 33'd466432104;
        test_addr[993] = 80;
        test_data[993] = 33'd3440150321;
        test_addr[994] = 81;
        test_data[994] = 33'd2609650108;
        test_addr[995] = 82;
        test_data[995] = 33'd5444661139;
        test_addr[996] = 83;
        test_data[996] = 33'd4471089093;
        test_addr[997] = 84;
        test_data[997] = 33'd389769389;
        test_addr[998] = 85;
        test_data[998] = 33'd7677719203;
        test_addr[999] = 86;
        test_data[999] = 33'd623629618;
        test_addr[1000] = 87;
        test_data[1000] = 33'd3303907992;
        test_addr[1001] = 88;
        test_data[1001] = 33'd8526148215;
        test_addr[1002] = 418;
        test_data[1002] = 33'd1591263160;
        test_addr[1003] = 420;
        test_data[1003] = 33'd443838194;
        test_addr[1004] = 421;
        test_data[1004] = 33'd3567358548;
        test_addr[1005] = 422;
        test_data[1005] = 33'd2973342047;
        test_addr[1006] = 423;
        test_data[1006] = 33'd1673945276;
        test_addr[1007] = 424;
        test_data[1007] = 33'd458707520;
        test_addr[1008] = 425;
        test_data[1008] = 33'd2344341674;
        test_addr[1009] = 426;
        test_data[1009] = 33'd5411200159;
        test_addr[1010] = 419;
        test_data[1010] = 33'd188335908;
        test_addr[1011] = 824;
        test_data[1011] = 33'd3204893334;
        test_addr[1012] = 420;
        test_data[1012] = 33'd5402362969;
        test_addr[1013] = 421;
        test_data[1013] = 33'd3567358548;
        test_addr[1014] = 422;
        test_data[1014] = 33'd7599357097;
        test_addr[1015] = 423;
        test_data[1015] = 33'd7245491000;
        test_addr[1016] = 424;
        test_data[1016] = 33'd458707520;
        test_addr[1017] = 425;
        test_data[1017] = 33'd2344341674;
        test_addr[1018] = 426;
        test_data[1018] = 33'd1116232863;
        test_addr[1019] = 427;
        test_data[1019] = 33'd1979928705;
        test_addr[1020] = 428;
        test_data[1020] = 33'd1479974522;
        test_addr[1021] = 429;
        test_data[1021] = 33'd3385333427;
        test_addr[1022] = 430;
        test_data[1022] = 33'd2489047385;
        test_addr[1023] = 431;
        test_data[1023] = 33'd5189287196;
        test_addr[1024] = 432;
        test_data[1024] = 33'd1474827311;
        test_addr[1025] = 638;
        test_data[1025] = 33'd881995127;
        test_addr[1026] = 639;
        test_data[1026] = 33'd1193599707;
        test_addr[1027] = 640;
        test_data[1027] = 33'd4856037743;
        test_addr[1028] = 641;
        test_data[1028] = 33'd2087204287;
        test_addr[1029] = 642;
        test_data[1029] = 33'd5066597340;
        test_addr[1030] = 643;
        test_data[1030] = 33'd8195005945;
        test_addr[1031] = 644;
        test_data[1031] = 33'd3175733827;
        test_addr[1032] = 645;
        test_data[1032] = 33'd2042867590;
        test_addr[1033] = 646;
        test_data[1033] = 33'd1737372841;
        test_addr[1034] = 647;
        test_data[1034] = 33'd3927182985;
        test_addr[1035] = 648;
        test_data[1035] = 33'd3673972943;
        test_addr[1036] = 649;
        test_data[1036] = 33'd2151483163;
        test_addr[1037] = 650;
        test_data[1037] = 33'd4155655242;
        test_addr[1038] = 433;
        test_data[1038] = 33'd7200177940;
        test_addr[1039] = 434;
        test_data[1039] = 33'd3881600915;
        test_addr[1040] = 435;
        test_data[1040] = 33'd1781223650;
        test_addr[1041] = 997;
        test_data[1041] = 33'd6740411736;
        test_addr[1042] = 998;
        test_data[1042] = 33'd5814685248;
        test_addr[1043] = 999;
        test_data[1043] = 33'd811944595;
        test_addr[1044] = 1000;
        test_data[1044] = 33'd5701976648;
        test_addr[1045] = 1001;
        test_data[1045] = 33'd3133226956;
        test_addr[1046] = 1002;
        test_data[1046] = 33'd1816079453;
        test_addr[1047] = 1003;
        test_data[1047] = 33'd4571456636;
        test_addr[1048] = 436;
        test_data[1048] = 33'd1024435444;
        test_addr[1049] = 437;
        test_data[1049] = 33'd390516077;
        test_addr[1050] = 438;
        test_data[1050] = 33'd3957892093;
        test_addr[1051] = 439;
        test_data[1051] = 33'd387768256;
        test_addr[1052] = 440;
        test_data[1052] = 33'd118271122;
        test_addr[1053] = 441;
        test_data[1053] = 33'd3910731565;
        test_addr[1054] = 442;
        test_data[1054] = 33'd4730441146;
        test_addr[1055] = 443;
        test_data[1055] = 33'd2309805798;
        test_addr[1056] = 444;
        test_data[1056] = 33'd4533997437;
        test_addr[1057] = 445;
        test_data[1057] = 33'd57979874;
        test_addr[1058] = 446;
        test_data[1058] = 33'd185249361;
        test_addr[1059] = 447;
        test_data[1059] = 33'd7785708212;
        test_addr[1060] = 448;
        test_data[1060] = 33'd4524420053;
        test_addr[1061] = 449;
        test_data[1061] = 33'd2000661367;
        test_addr[1062] = 450;
        test_data[1062] = 33'd1220832376;
        test_addr[1063] = 451;
        test_data[1063] = 33'd2278524113;
        test_addr[1064] = 452;
        test_data[1064] = 33'd4472183568;
        test_addr[1065] = 453;
        test_data[1065] = 33'd2615425596;
        test_addr[1066] = 454;
        test_data[1066] = 33'd6567695374;
        test_addr[1067] = 455;
        test_data[1067] = 33'd5912745263;
        test_addr[1068] = 456;
        test_data[1068] = 33'd1297742875;
        test_addr[1069] = 654;
        test_data[1069] = 33'd5725808381;
        test_addr[1070] = 655;
        test_data[1070] = 33'd1564587862;
        test_addr[1071] = 656;
        test_data[1071] = 33'd1587342591;
        test_addr[1072] = 657;
        test_data[1072] = 33'd2971496127;
        test_addr[1073] = 658;
        test_data[1073] = 33'd6300500720;
        test_addr[1074] = 659;
        test_data[1074] = 33'd4171986551;
        test_addr[1075] = 660;
        test_data[1075] = 33'd3089242911;
        test_addr[1076] = 661;
        test_data[1076] = 33'd507482648;
        test_addr[1077] = 662;
        test_data[1077] = 33'd8233406385;
        test_addr[1078] = 663;
        test_data[1078] = 33'd2975358863;
        test_addr[1079] = 664;
        test_data[1079] = 33'd7661659957;
        test_addr[1080] = 665;
        test_data[1080] = 33'd6625012026;
        test_addr[1081] = 666;
        test_data[1081] = 33'd3229102402;
        test_addr[1082] = 667;
        test_data[1082] = 33'd2248979690;
        test_addr[1083] = 668;
        test_data[1083] = 33'd2810872159;
        test_addr[1084] = 669;
        test_data[1084] = 33'd7146106679;
        test_addr[1085] = 457;
        test_data[1085] = 33'd2700525639;
        test_addr[1086] = 458;
        test_data[1086] = 33'd1845881788;
        test_addr[1087] = 459;
        test_data[1087] = 33'd582707416;
        test_addr[1088] = 460;
        test_data[1088] = 33'd3277373807;
        test_addr[1089] = 461;
        test_data[1089] = 33'd4878573432;
        test_addr[1090] = 488;
        test_data[1090] = 33'd8004619445;
        test_addr[1091] = 489;
        test_data[1091] = 33'd7113195223;
        test_addr[1092] = 462;
        test_data[1092] = 33'd8067760642;
        test_addr[1093] = 463;
        test_data[1093] = 33'd5569735010;
        test_addr[1094] = 464;
        test_data[1094] = 33'd1701612275;
        test_addr[1095] = 465;
        test_data[1095] = 33'd2952264133;
        test_addr[1096] = 466;
        test_data[1096] = 33'd2807963646;
        test_addr[1097] = 467;
        test_data[1097] = 33'd962725890;
        test_addr[1098] = 468;
        test_data[1098] = 33'd7168246071;
        test_addr[1099] = 469;
        test_data[1099] = 33'd1191579314;
        test_addr[1100] = 470;
        test_data[1100] = 33'd1183712898;
        test_addr[1101] = 775;
        test_data[1101] = 33'd4171009354;
        test_addr[1102] = 776;
        test_data[1102] = 33'd3596983855;
        test_addr[1103] = 777;
        test_data[1103] = 33'd3617657151;
        test_addr[1104] = 778;
        test_data[1104] = 33'd1257411684;
        test_addr[1105] = 779;
        test_data[1105] = 33'd8273649709;
        test_addr[1106] = 780;
        test_data[1106] = 33'd1167957788;
        test_addr[1107] = 781;
        test_data[1107] = 33'd5423482006;
        test_addr[1108] = 782;
        test_data[1108] = 33'd6947357753;
        test_addr[1109] = 783;
        test_data[1109] = 33'd7140426857;
        test_addr[1110] = 784;
        test_data[1110] = 33'd7660476717;
        test_addr[1111] = 785;
        test_data[1111] = 33'd8586299103;
        test_addr[1112] = 786;
        test_data[1112] = 33'd7990484284;
        test_addr[1113] = 787;
        test_data[1113] = 33'd5123258959;
        test_addr[1114] = 788;
        test_data[1114] = 33'd1105670773;
        test_addr[1115] = 789;
        test_data[1115] = 33'd911008138;
        test_addr[1116] = 471;
        test_data[1116] = 33'd7942050822;
        test_addr[1117] = 472;
        test_data[1117] = 33'd6439358734;
        test_addr[1118] = 473;
        test_data[1118] = 33'd2376303146;
        test_addr[1119] = 474;
        test_data[1119] = 33'd107046119;
        test_addr[1120] = 475;
        test_data[1120] = 33'd1588844006;
        test_addr[1121] = 476;
        test_data[1121] = 33'd5274340300;
        test_addr[1122] = 950;
        test_data[1122] = 33'd2459752245;
        test_addr[1123] = 951;
        test_data[1123] = 33'd3631193825;
        test_addr[1124] = 952;
        test_data[1124] = 33'd1791314849;
        test_addr[1125] = 953;
        test_data[1125] = 33'd2693867941;
        test_addr[1126] = 477;
        test_data[1126] = 33'd702771066;
        test_addr[1127] = 478;
        test_data[1127] = 33'd3853924173;
        test_addr[1128] = 54;
        test_data[1128] = 33'd7283787228;
        test_addr[1129] = 55;
        test_data[1129] = 33'd6525576188;
        test_addr[1130] = 56;
        test_data[1130] = 33'd5804565453;
        test_addr[1131] = 57;
        test_data[1131] = 33'd22011062;
        test_addr[1132] = 58;
        test_data[1132] = 33'd3203147784;
        test_addr[1133] = 59;
        test_data[1133] = 33'd1487397129;
        test_addr[1134] = 60;
        test_data[1134] = 33'd4664823303;
        test_addr[1135] = 61;
        test_data[1135] = 33'd2209095858;
        test_addr[1136] = 62;
        test_data[1136] = 33'd504570280;
        test_addr[1137] = 63;
        test_data[1137] = 33'd8438126187;
        test_addr[1138] = 64;
        test_data[1138] = 33'd6000401759;
        test_addr[1139] = 65;
        test_data[1139] = 33'd4169485515;
        test_addr[1140] = 66;
        test_data[1140] = 33'd3795061744;
        test_addr[1141] = 67;
        test_data[1141] = 33'd2781999553;
        test_addr[1142] = 68;
        test_data[1142] = 33'd2440392340;
        test_addr[1143] = 69;
        test_data[1143] = 33'd7284517722;
        test_addr[1144] = 70;
        test_data[1144] = 33'd3874690545;
        test_addr[1145] = 71;
        test_data[1145] = 33'd1800624896;
        test_addr[1146] = 72;
        test_data[1146] = 33'd3745474962;
        test_addr[1147] = 73;
        test_data[1147] = 33'd7724627947;
        test_addr[1148] = 74;
        test_data[1148] = 33'd1195861608;
        test_addr[1149] = 75;
        test_data[1149] = 33'd7685967673;
        test_addr[1150] = 76;
        test_data[1150] = 33'd1051232611;
        test_addr[1151] = 77;
        test_data[1151] = 33'd6717808536;
        test_addr[1152] = 78;
        test_data[1152] = 33'd3591490314;
        test_addr[1153] = 479;
        test_data[1153] = 33'd2750306313;
        test_addr[1154] = 480;
        test_data[1154] = 33'd1372344996;
        test_addr[1155] = 481;
        test_data[1155] = 33'd7289728586;
        test_addr[1156] = 482;
        test_data[1156] = 33'd2222178533;
        test_addr[1157] = 483;
        test_data[1157] = 33'd3017205182;
        test_addr[1158] = 484;
        test_data[1158] = 33'd1185966804;
        test_addr[1159] = 10;
        test_data[1159] = 33'd4271687727;
        test_addr[1160] = 11;
        test_data[1160] = 33'd3967754806;
        test_addr[1161] = 12;
        test_data[1161] = 33'd1768449257;
        test_addr[1162] = 13;
        test_data[1162] = 33'd716472127;
        test_addr[1163] = 14;
        test_data[1163] = 33'd6926169710;
        test_addr[1164] = 485;
        test_data[1164] = 33'd6077775508;
        test_addr[1165] = 486;
        test_data[1165] = 33'd2334539005;
        test_addr[1166] = 487;
        test_data[1166] = 33'd3597154848;
        test_addr[1167] = 488;
        test_data[1167] = 33'd3709652149;
        test_addr[1168] = 219;
        test_data[1168] = 33'd3593970920;
        test_addr[1169] = 220;
        test_data[1169] = 33'd5023328405;
        test_addr[1170] = 221;
        test_data[1170] = 33'd6652082891;
        test_addr[1171] = 222;
        test_data[1171] = 33'd4233733742;
        test_addr[1172] = 223;
        test_data[1172] = 33'd308136402;
        test_addr[1173] = 224;
        test_data[1173] = 33'd7627397883;
        test_addr[1174] = 225;
        test_data[1174] = 33'd1255812106;
        test_addr[1175] = 226;
        test_data[1175] = 33'd7178749101;
        test_addr[1176] = 227;
        test_data[1176] = 33'd4650952586;
        test_addr[1177] = 228;
        test_data[1177] = 33'd2819019937;
        test_addr[1178] = 229;
        test_data[1178] = 33'd845232644;
        test_addr[1179] = 230;
        test_data[1179] = 33'd92067608;
        test_addr[1180] = 231;
        test_data[1180] = 33'd4459237376;
        test_addr[1181] = 232;
        test_data[1181] = 33'd4110523392;
        test_addr[1182] = 233;
        test_data[1182] = 33'd6599594934;
        test_addr[1183] = 234;
        test_data[1183] = 33'd7847118232;
        test_addr[1184] = 235;
        test_data[1184] = 33'd1995153683;
        test_addr[1185] = 489;
        test_data[1185] = 33'd2818227927;
        test_addr[1186] = 490;
        test_data[1186] = 33'd541064026;
        test_addr[1187] = 491;
        test_data[1187] = 33'd4919423175;
        test_addr[1188] = 492;
        test_data[1188] = 33'd5468665486;
        test_addr[1189] = 493;
        test_data[1189] = 33'd1126176295;
        test_addr[1190] = 494;
        test_data[1190] = 33'd2546758818;
        test_addr[1191] = 495;
        test_data[1191] = 33'd1266991624;
        test_addr[1192] = 496;
        test_data[1192] = 33'd4987737681;
        test_addr[1193] = 497;
        test_data[1193] = 33'd4946439286;
        test_addr[1194] = 498;
        test_data[1194] = 33'd1319694326;
        test_addr[1195] = 853;
        test_data[1195] = 33'd782842199;
        test_addr[1196] = 854;
        test_data[1196] = 33'd4381862831;
        test_addr[1197] = 855;
        test_data[1197] = 33'd3155227187;
        test_addr[1198] = 856;
        test_data[1198] = 33'd7030537960;
        test_addr[1199] = 499;
        test_data[1199] = 33'd2620324755;
        test_addr[1200] = 500;
        test_data[1200] = 33'd1324133867;
        test_addr[1201] = 501;
        test_data[1201] = 33'd2750530624;
        test_addr[1202] = 502;
        test_data[1202] = 33'd8148991678;
        test_addr[1203] = 503;
        test_data[1203] = 33'd5138690788;
        test_addr[1204] = 504;
        test_data[1204] = 33'd951027809;
        test_addr[1205] = 505;
        test_data[1205] = 33'd1706057765;
        test_addr[1206] = 506;
        test_data[1206] = 33'd5142876609;
        test_addr[1207] = 507;
        test_data[1207] = 33'd8101750497;
        test_addr[1208] = 508;
        test_data[1208] = 33'd3779675938;
        test_addr[1209] = 509;
        test_data[1209] = 33'd1248057624;
        test_addr[1210] = 510;
        test_data[1210] = 33'd7367678905;
        test_addr[1211] = 511;
        test_data[1211] = 33'd3342970419;
        test_addr[1212] = 512;
        test_data[1212] = 33'd283576485;
        test_addr[1213] = 513;
        test_data[1213] = 33'd3832833658;
        test_addr[1214] = 514;
        test_data[1214] = 33'd6036200334;
        test_addr[1215] = 515;
        test_data[1215] = 33'd4175963926;
        test_addr[1216] = 516;
        test_data[1216] = 33'd7226984075;
        test_addr[1217] = 517;
        test_data[1217] = 33'd1173365637;
        test_addr[1218] = 518;
        test_data[1218] = 33'd2424591448;
        test_addr[1219] = 519;
        test_data[1219] = 33'd2472061153;
        test_addr[1220] = 520;
        test_data[1220] = 33'd2499178703;
        test_addr[1221] = 521;
        test_data[1221] = 33'd8240402564;
        test_addr[1222] = 522;
        test_data[1222] = 33'd2119484876;
        test_addr[1223] = 523;
        test_data[1223] = 33'd2084861691;
        test_addr[1224] = 524;
        test_data[1224] = 33'd4169713201;
        test_addr[1225] = 525;
        test_data[1225] = 33'd2372613957;
        test_addr[1226] = 526;
        test_data[1226] = 33'd5175506030;
        test_addr[1227] = 527;
        test_data[1227] = 33'd1738182943;
        test_addr[1228] = 528;
        test_data[1228] = 33'd4959772114;
        test_addr[1229] = 529;
        test_data[1229] = 33'd6903503381;
        test_addr[1230] = 530;
        test_data[1230] = 33'd1199134247;
        test_addr[1231] = 531;
        test_data[1231] = 33'd5340479159;
        test_addr[1232] = 532;
        test_data[1232] = 33'd1098075619;
        test_addr[1233] = 533;
        test_data[1233] = 33'd5115261679;
        test_addr[1234] = 534;
        test_data[1234] = 33'd627486554;
        test_addr[1235] = 535;
        test_data[1235] = 33'd2501250615;
        test_addr[1236] = 536;
        test_data[1236] = 33'd4241396361;
        test_addr[1237] = 537;
        test_data[1237] = 33'd1845215902;
        test_addr[1238] = 172;
        test_data[1238] = 33'd8492972273;
        test_addr[1239] = 173;
        test_data[1239] = 33'd5999007414;
        test_addr[1240] = 174;
        test_data[1240] = 33'd6580079718;
        test_addr[1241] = 175;
        test_data[1241] = 33'd3567745488;
        test_addr[1242] = 176;
        test_data[1242] = 33'd6717825895;
        test_addr[1243] = 177;
        test_data[1243] = 33'd2295881178;
        test_addr[1244] = 178;
        test_data[1244] = 33'd5040266672;
        test_addr[1245] = 179;
        test_data[1245] = 33'd2886227464;
        test_addr[1246] = 180;
        test_data[1246] = 33'd4240384840;
        test_addr[1247] = 181;
        test_data[1247] = 33'd6451215601;
        test_addr[1248] = 182;
        test_data[1248] = 33'd1222529405;
        test_addr[1249] = 183;
        test_data[1249] = 33'd4192569996;
        test_addr[1250] = 184;
        test_data[1250] = 33'd961772350;
        test_addr[1251] = 185;
        test_data[1251] = 33'd3717107221;
        test_addr[1252] = 186;
        test_data[1252] = 33'd2175561490;
        test_addr[1253] = 187;
        test_data[1253] = 33'd3131077888;
        test_addr[1254] = 188;
        test_data[1254] = 33'd128496091;
        test_addr[1255] = 189;
        test_data[1255] = 33'd133639369;
        test_addr[1256] = 190;
        test_data[1256] = 33'd4284820396;
        test_addr[1257] = 191;
        test_data[1257] = 33'd3150765077;
        test_addr[1258] = 192;
        test_data[1258] = 33'd275041321;
        test_addr[1259] = 193;
        test_data[1259] = 33'd122598896;
        test_addr[1260] = 194;
        test_data[1260] = 33'd8335297207;
        test_addr[1261] = 195;
        test_data[1261] = 33'd3241511229;
        test_addr[1262] = 196;
        test_data[1262] = 33'd1811402878;
        test_addr[1263] = 197;
        test_data[1263] = 33'd5455018927;
        test_addr[1264] = 198;
        test_data[1264] = 33'd1771443269;
        test_addr[1265] = 199;
        test_data[1265] = 33'd4580577277;
        test_addr[1266] = 200;
        test_data[1266] = 33'd6602403768;
        test_addr[1267] = 201;
        test_data[1267] = 33'd1922645171;
        test_addr[1268] = 202;
        test_data[1268] = 33'd5219335820;
        test_addr[1269] = 203;
        test_data[1269] = 33'd1663091370;
        test_addr[1270] = 204;
        test_data[1270] = 33'd7368337612;
        test_addr[1271] = 538;
        test_data[1271] = 33'd2288013246;
        test_addr[1272] = 539;
        test_data[1272] = 33'd2749828337;
        test_addr[1273] = 540;
        test_data[1273] = 33'd30470061;
        test_addr[1274] = 541;
        test_data[1274] = 33'd2310349212;
        test_addr[1275] = 542;
        test_data[1275] = 33'd2967622748;
        test_addr[1276] = 543;
        test_data[1276] = 33'd4593646050;
        test_addr[1277] = 544;
        test_data[1277] = 33'd3477380391;
        test_addr[1278] = 545;
        test_data[1278] = 33'd5924966091;
        test_addr[1279] = 546;
        test_data[1279] = 33'd8109295558;
        test_addr[1280] = 547;
        test_data[1280] = 33'd3210837133;
        test_addr[1281] = 548;
        test_data[1281] = 33'd1180199925;
        test_addr[1282] = 549;
        test_data[1282] = 33'd6772317964;
        test_addr[1283] = 550;
        test_data[1283] = 33'd2009710279;
        test_addr[1284] = 551;
        test_data[1284] = 33'd318746959;
        test_addr[1285] = 552;
        test_data[1285] = 33'd6523742868;
        test_addr[1286] = 387;
        test_data[1286] = 33'd3152915513;
        test_addr[1287] = 388;
        test_data[1287] = 33'd2217298716;
        test_addr[1288] = 389;
        test_data[1288] = 33'd2233888802;
        test_addr[1289] = 390;
        test_data[1289] = 33'd3947964093;
        test_addr[1290] = 391;
        test_data[1290] = 33'd4156755592;
        test_addr[1291] = 392;
        test_data[1291] = 33'd4621624781;
        test_addr[1292] = 393;
        test_data[1292] = 33'd3584816215;
        test_addr[1293] = 394;
        test_data[1293] = 33'd6638130426;
        test_addr[1294] = 395;
        test_data[1294] = 33'd7844710652;
        test_addr[1295] = 396;
        test_data[1295] = 33'd179786261;
        test_addr[1296] = 397;
        test_data[1296] = 33'd8169636037;
        test_addr[1297] = 553;
        test_data[1297] = 33'd298968730;
        test_addr[1298] = 554;
        test_data[1298] = 33'd3262924390;
        test_addr[1299] = 555;
        test_data[1299] = 33'd449821878;
        test_addr[1300] = 556;
        test_data[1300] = 33'd2994603037;
        test_addr[1301] = 557;
        test_data[1301] = 33'd2415573794;
        test_addr[1302] = 558;
        test_data[1302] = 33'd3010760443;
        test_addr[1303] = 559;
        test_data[1303] = 33'd455792188;
        test_addr[1304] = 560;
        test_data[1304] = 33'd6599501376;
        test_addr[1305] = 561;
        test_data[1305] = 33'd1362019700;
        test_addr[1306] = 56;
        test_data[1306] = 33'd8485920423;
        test_addr[1307] = 57;
        test_data[1307] = 33'd6615721998;
        test_addr[1308] = 58;
        test_data[1308] = 33'd3203147784;
        test_addr[1309] = 562;
        test_data[1309] = 33'd286708441;
        test_addr[1310] = 563;
        test_data[1310] = 33'd38688635;
        test_addr[1311] = 564;
        test_data[1311] = 33'd2631069284;
        test_addr[1312] = 565;
        test_data[1312] = 33'd6498517760;
        test_addr[1313] = 566;
        test_data[1313] = 33'd3270728084;
        test_addr[1314] = 567;
        test_data[1314] = 33'd5124711129;
        test_addr[1315] = 568;
        test_data[1315] = 33'd352858729;
        test_addr[1316] = 569;
        test_data[1316] = 33'd1734513920;
        test_addr[1317] = 570;
        test_data[1317] = 33'd5312316431;
        test_addr[1318] = 898;
        test_data[1318] = 33'd6070265227;
        test_addr[1319] = 899;
        test_data[1319] = 33'd4140880084;
        test_addr[1320] = 900;
        test_data[1320] = 33'd6376673680;
        test_addr[1321] = 901;
        test_data[1321] = 33'd5899833155;
        test_addr[1322] = 902;
        test_data[1322] = 33'd3561446271;
        test_addr[1323] = 571;
        test_data[1323] = 33'd2564920536;
        test_addr[1324] = 572;
        test_data[1324] = 33'd2320974549;
        test_addr[1325] = 197;
        test_data[1325] = 33'd1160051631;
        test_addr[1326] = 198;
        test_data[1326] = 33'd1771443269;
        test_addr[1327] = 199;
        test_data[1327] = 33'd285609981;
        test_addr[1328] = 200;
        test_data[1328] = 33'd5916701174;
        test_addr[1329] = 201;
        test_data[1329] = 33'd7419932114;
        test_addr[1330] = 202;
        test_data[1330] = 33'd8499463203;
        test_addr[1331] = 203;
        test_data[1331] = 33'd1663091370;
        test_addr[1332] = 204;
        test_data[1332] = 33'd3073370316;
        test_addr[1333] = 205;
        test_data[1333] = 33'd349509858;
        test_addr[1334] = 206;
        test_data[1334] = 33'd871555750;
        test_addr[1335] = 207;
        test_data[1335] = 33'd3823761644;
        test_addr[1336] = 208;
        test_data[1336] = 33'd3010632164;
        test_addr[1337] = 209;
        test_data[1337] = 33'd2101436476;
        test_addr[1338] = 210;
        test_data[1338] = 33'd4686413679;
        test_addr[1339] = 211;
        test_data[1339] = 33'd3337632621;
        test_addr[1340] = 212;
        test_data[1340] = 33'd2977847200;
        test_addr[1341] = 213;
        test_data[1341] = 33'd371999850;
        test_addr[1342] = 214;
        test_data[1342] = 33'd5262987318;
        test_addr[1343] = 215;
        test_data[1343] = 33'd2179149214;
        test_addr[1344] = 216;
        test_data[1344] = 33'd5003308831;
        test_addr[1345] = 217;
        test_data[1345] = 33'd797224449;
        test_addr[1346] = 218;
        test_data[1346] = 33'd5477752146;
        test_addr[1347] = 219;
        test_data[1347] = 33'd6984031259;
        test_addr[1348] = 220;
        test_data[1348] = 33'd728361109;
        test_addr[1349] = 221;
        test_data[1349] = 33'd6074992176;
        test_addr[1350] = 222;
        test_data[1350] = 33'd4233733742;
        test_addr[1351] = 223;
        test_data[1351] = 33'd8065317518;
        test_addr[1352] = 224;
        test_data[1352] = 33'd3332430587;
        test_addr[1353] = 225;
        test_data[1353] = 33'd4501064444;
        test_addr[1354] = 226;
        test_data[1354] = 33'd2883781805;
        test_addr[1355] = 227;
        test_data[1355] = 33'd355985290;
        test_addr[1356] = 228;
        test_data[1356] = 33'd2819019937;
        test_addr[1357] = 229;
        test_data[1357] = 33'd845232644;
        test_addr[1358] = 230;
        test_data[1358] = 33'd7707061078;
        test_addr[1359] = 231;
        test_data[1359] = 33'd164270080;
        test_addr[1360] = 232;
        test_data[1360] = 33'd4406171327;
        test_addr[1361] = 233;
        test_data[1361] = 33'd2304627638;
        test_addr[1362] = 234;
        test_data[1362] = 33'd3552150936;
        test_addr[1363] = 235;
        test_data[1363] = 33'd1995153683;
        test_addr[1364] = 236;
        test_data[1364] = 33'd3308823479;
        test_addr[1365] = 237;
        test_data[1365] = 33'd7583394011;
        test_addr[1366] = 238;
        test_data[1366] = 33'd6050016741;
        test_addr[1367] = 573;
        test_data[1367] = 33'd4530893709;
        test_addr[1368] = 574;
        test_data[1368] = 33'd1311509596;
        test_addr[1369] = 575;
        test_data[1369] = 33'd1340627649;
        test_addr[1370] = 576;
        test_data[1370] = 33'd2352940238;
        test_addr[1371] = 577;
        test_data[1371] = 33'd6088920071;
        test_addr[1372] = 578;
        test_data[1372] = 33'd7491261717;
        test_addr[1373] = 579;
        test_data[1373] = 33'd1094013198;
        test_addr[1374] = 580;
        test_data[1374] = 33'd1233267658;
        test_addr[1375] = 581;
        test_data[1375] = 33'd962066425;
        test_addr[1376] = 582;
        test_data[1376] = 33'd3179541911;
        test_addr[1377] = 583;
        test_data[1377] = 33'd2231704842;
        test_addr[1378] = 584;
        test_data[1378] = 33'd1490217735;
        test_addr[1379] = 585;
        test_data[1379] = 33'd1270660057;
        test_addr[1380] = 586;
        test_data[1380] = 33'd1844798620;
        test_addr[1381] = 587;
        test_data[1381] = 33'd6304397302;
        test_addr[1382] = 588;
        test_data[1382] = 33'd1893529001;
        test_addr[1383] = 589;
        test_data[1383] = 33'd3514985912;
        test_addr[1384] = 590;
        test_data[1384] = 33'd2083229337;
        test_addr[1385] = 591;
        test_data[1385] = 33'd4798286920;
        test_addr[1386] = 592;
        test_data[1386] = 33'd1467139886;
        test_addr[1387] = 593;
        test_data[1387] = 33'd704520665;
        test_addr[1388] = 594;
        test_data[1388] = 33'd499927349;
        test_addr[1389] = 595;
        test_data[1389] = 33'd2612499855;
        test_addr[1390] = 596;
        test_data[1390] = 33'd2164998835;
        test_addr[1391] = 597;
        test_data[1391] = 33'd8564079049;
        test_addr[1392] = 598;
        test_data[1392] = 33'd3698561184;
        test_addr[1393] = 599;
        test_data[1393] = 33'd2621666958;
        test_addr[1394] = 600;
        test_data[1394] = 33'd5324017021;
        test_addr[1395] = 601;
        test_data[1395] = 33'd647592843;
        test_addr[1396] = 602;
        test_data[1396] = 33'd1224924786;
        test_addr[1397] = 603;
        test_data[1397] = 33'd6342231797;
        test_addr[1398] = 604;
        test_data[1398] = 33'd152904658;
        test_addr[1399] = 256;
        test_data[1399] = 33'd7648588057;
        test_addr[1400] = 605;
        test_data[1400] = 33'd4068052147;
        test_addr[1401] = 606;
        test_data[1401] = 33'd906696308;
        test_addr[1402] = 607;
        test_data[1402] = 33'd6382266354;
        test_addr[1403] = 608;
        test_data[1403] = 33'd3635138265;
        test_addr[1404] = 609;
        test_data[1404] = 33'd6437018279;
        test_addr[1405] = 610;
        test_data[1405] = 33'd2988230185;
        test_addr[1406] = 611;
        test_data[1406] = 33'd180393329;
        test_addr[1407] = 612;
        test_data[1407] = 33'd2469017315;
        test_addr[1408] = 613;
        test_data[1408] = 33'd3646976116;
        test_addr[1409] = 614;
        test_data[1409] = 33'd7923231515;
        test_addr[1410] = 615;
        test_data[1410] = 33'd995474728;
        test_addr[1411] = 616;
        test_data[1411] = 33'd1306428470;
        test_addr[1412] = 617;
        test_data[1412] = 33'd5726785392;
        test_addr[1413] = 308;
        test_data[1413] = 33'd2611705428;
        test_addr[1414] = 309;
        test_data[1414] = 33'd3941608837;
        test_addr[1415] = 618;
        test_data[1415] = 33'd7439529767;
        test_addr[1416] = 619;
        test_data[1416] = 33'd4949805919;
        test_addr[1417] = 620;
        test_data[1417] = 33'd5456429013;
        test_addr[1418] = 621;
        test_data[1418] = 33'd723470077;
        test_addr[1419] = 622;
        test_data[1419] = 33'd6937931629;
        test_addr[1420] = 623;
        test_data[1420] = 33'd2813751329;
        test_addr[1421] = 624;
        test_data[1421] = 33'd2812841878;
        test_addr[1422] = 625;
        test_data[1422] = 33'd2462103418;
        test_addr[1423] = 626;
        test_data[1423] = 33'd7982824441;
        test_addr[1424] = 627;
        test_data[1424] = 33'd5545982797;
        test_addr[1425] = 628;
        test_data[1425] = 33'd2469942537;
        test_addr[1426] = 629;
        test_data[1426] = 33'd3332408304;
        test_addr[1427] = 630;
        test_data[1427] = 33'd4675669049;
        test_addr[1428] = 631;
        test_data[1428] = 33'd7554920012;
        test_addr[1429] = 632;
        test_data[1429] = 33'd3201343516;
        test_addr[1430] = 846;
        test_data[1430] = 33'd3157279990;
        test_addr[1431] = 847;
        test_data[1431] = 33'd4178636307;
        test_addr[1432] = 633;
        test_data[1432] = 33'd1874676766;
        test_addr[1433] = 634;
        test_data[1433] = 33'd954992338;
        test_addr[1434] = 635;
        test_data[1434] = 33'd8269660053;
        test_addr[1435] = 636;
        test_data[1435] = 33'd4218479966;
        test_addr[1436] = 637;
        test_data[1436] = 33'd3795165725;
        test_addr[1437] = 638;
        test_data[1437] = 33'd881995127;
        test_addr[1438] = 639;
        test_data[1438] = 33'd6545300217;
        test_addr[1439] = 640;
        test_data[1439] = 33'd561070447;
        test_addr[1440] = 641;
        test_data[1440] = 33'd2087204287;
        test_addr[1441] = 745;
        test_data[1441] = 33'd5627963735;
        test_addr[1442] = 746;
        test_data[1442] = 33'd5551477754;
        test_addr[1443] = 747;
        test_data[1443] = 33'd6515224038;
        test_addr[1444] = 748;
        test_data[1444] = 33'd1521829790;
        test_addr[1445] = 749;
        test_data[1445] = 33'd8247155540;
        test_addr[1446] = 750;
        test_data[1446] = 33'd282558174;
        test_addr[1447] = 642;
        test_data[1447] = 33'd771630044;
        test_addr[1448] = 643;
        test_data[1448] = 33'd3900038649;
        test_addr[1449] = 644;
        test_data[1449] = 33'd3175733827;
        test_addr[1450] = 645;
        test_data[1450] = 33'd8364755595;
        test_addr[1451] = 646;
        test_data[1451] = 33'd1737372841;
        test_addr[1452] = 647;
        test_data[1452] = 33'd5785972390;
        test_addr[1453] = 648;
        test_data[1453] = 33'd6525490539;
        test_addr[1454] = 649;
        test_data[1454] = 33'd7052366868;
        test_addr[1455] = 650;
        test_data[1455] = 33'd7328578652;
        test_addr[1456] = 651;
        test_data[1456] = 33'd2006915388;
        test_addr[1457] = 652;
        test_data[1457] = 33'd3998291136;
        test_addr[1458] = 653;
        test_data[1458] = 33'd5236861111;
        test_addr[1459] = 654;
        test_data[1459] = 33'd1430841085;
        test_addr[1460] = 655;
        test_data[1460] = 33'd1564587862;
        test_addr[1461] = 656;
        test_data[1461] = 33'd1587342591;
        test_addr[1462] = 657;
        test_data[1462] = 33'd2971496127;
        test_addr[1463] = 658;
        test_data[1463] = 33'd7897220974;
        test_addr[1464] = 659;
        test_data[1464] = 33'd5708950281;
        test_addr[1465] = 660;
        test_data[1465] = 33'd3089242911;
        test_addr[1466] = 661;
        test_data[1466] = 33'd507482648;
        test_addr[1467] = 662;
        test_data[1467] = 33'd3938439089;
        test_addr[1468] = 663;
        test_data[1468] = 33'd6696485811;
        test_addr[1469] = 334;
        test_data[1469] = 33'd4662372669;
        test_addr[1470] = 335;
        test_data[1470] = 33'd6465099796;
        test_addr[1471] = 336;
        test_data[1471] = 33'd2188727585;
        test_addr[1472] = 337;
        test_data[1472] = 33'd7333966563;
        test_addr[1473] = 338;
        test_data[1473] = 33'd5195610624;
        test_addr[1474] = 339;
        test_data[1474] = 33'd2387661980;
        test_addr[1475] = 340;
        test_data[1475] = 33'd451413948;
        test_addr[1476] = 341;
        test_data[1476] = 33'd6269461644;
        test_addr[1477] = 664;
        test_data[1477] = 33'd3366692661;
        test_addr[1478] = 665;
        test_data[1478] = 33'd2330044730;
        test_addr[1479] = 53;
        test_data[1479] = 33'd6392110754;
        test_addr[1480] = 54;
        test_data[1480] = 33'd2988819932;
        test_addr[1481] = 55;
        test_data[1481] = 33'd2230608892;
        test_addr[1482] = 56;
        test_data[1482] = 33'd4190953127;
        test_addr[1483] = 57;
        test_data[1483] = 33'd2320754702;
        test_addr[1484] = 58;
        test_data[1484] = 33'd3203147784;
        test_addr[1485] = 59;
        test_data[1485] = 33'd7712740041;
        test_addr[1486] = 60;
        test_data[1486] = 33'd6125236980;
        test_addr[1487] = 61;
        test_data[1487] = 33'd2209095858;
        test_addr[1488] = 666;
        test_data[1488] = 33'd4923885202;
        test_addr[1489] = 667;
        test_data[1489] = 33'd7929291799;
        test_addr[1490] = 668;
        test_data[1490] = 33'd2810872159;
        test_addr[1491] = 669;
        test_data[1491] = 33'd4395709248;
        test_addr[1492] = 976;
        test_data[1492] = 33'd888555328;
        test_addr[1493] = 977;
        test_data[1493] = 33'd871000283;
        test_addr[1494] = 978;
        test_data[1494] = 33'd5862497060;
        test_addr[1495] = 979;
        test_data[1495] = 33'd3552257411;
        test_addr[1496] = 980;
        test_data[1496] = 33'd3721886817;
        test_addr[1497] = 981;
        test_data[1497] = 33'd4461748535;
        test_addr[1498] = 982;
        test_data[1498] = 33'd2064422908;
        test_addr[1499] = 983;
        test_data[1499] = 33'd6933935485;
        test_addr[1500] = 984;
        test_data[1500] = 33'd447706912;
        test_addr[1501] = 985;
        test_data[1501] = 33'd3871310064;
        test_addr[1502] = 986;
        test_data[1502] = 33'd2041805604;
        test_addr[1503] = 987;
        test_data[1503] = 33'd730636411;
        test_addr[1504] = 988;
        test_data[1504] = 33'd1189533474;
        test_addr[1505] = 989;
        test_data[1505] = 33'd5953280263;
        test_addr[1506] = 990;
        test_data[1506] = 33'd431413773;
        test_addr[1507] = 670;
        test_data[1507] = 33'd3197879796;
        test_addr[1508] = 671;
        test_data[1508] = 33'd3754236325;
        test_addr[1509] = 672;
        test_data[1509] = 33'd1411628437;
        test_addr[1510] = 673;
        test_data[1510] = 33'd1252547980;
        test_addr[1511] = 674;
        test_data[1511] = 33'd5383586391;
        test_addr[1512] = 675;
        test_data[1512] = 33'd3065041083;
        test_addr[1513] = 676;
        test_data[1513] = 33'd2458873297;
        test_addr[1514] = 677;
        test_data[1514] = 33'd3780631796;
        test_addr[1515] = 678;
        test_data[1515] = 33'd2431021203;
        test_addr[1516] = 679;
        test_data[1516] = 33'd2933532045;
        test_addr[1517] = 600;
        test_data[1517] = 33'd1029049725;
        test_addr[1518] = 601;
        test_data[1518] = 33'd647592843;
        test_addr[1519] = 602;
        test_data[1519] = 33'd1224924786;
        test_addr[1520] = 603;
        test_data[1520] = 33'd7860453720;
        test_addr[1521] = 604;
        test_data[1521] = 33'd6120391020;
        test_addr[1522] = 680;
        test_data[1522] = 33'd1881433713;
        test_addr[1523] = 681;
        test_data[1523] = 33'd1760731286;
        test_addr[1524] = 682;
        test_data[1524] = 33'd3793810237;
        test_addr[1525] = 683;
        test_data[1525] = 33'd1205808495;
        test_addr[1526] = 684;
        test_data[1526] = 33'd4251338616;
        test_addr[1527] = 685;
        test_data[1527] = 33'd1848469040;
        test_addr[1528] = 686;
        test_data[1528] = 33'd3756581141;
        test_addr[1529] = 687;
        test_data[1529] = 33'd5272397510;
        test_addr[1530] = 688;
        test_data[1530] = 33'd3658468012;
        test_addr[1531] = 689;
        test_data[1531] = 33'd1050422211;
        test_addr[1532] = 690;
        test_data[1532] = 33'd7271430356;
        test_addr[1533] = 691;
        test_data[1533] = 33'd1533424138;
        test_addr[1534] = 692;
        test_data[1534] = 33'd1185532734;
        test_addr[1535] = 693;
        test_data[1535] = 33'd1966776275;
        test_addr[1536] = 453;
        test_data[1536] = 33'd2615425596;
        test_addr[1537] = 454;
        test_data[1537] = 33'd2272728078;
        test_addr[1538] = 455;
        test_data[1538] = 33'd7345893899;
        test_addr[1539] = 456;
        test_data[1539] = 33'd1297742875;
        test_addr[1540] = 457;
        test_data[1540] = 33'd2700525639;
        test_addr[1541] = 458;
        test_data[1541] = 33'd6991938668;
        test_addr[1542] = 459;
        test_data[1542] = 33'd582707416;
        test_addr[1543] = 460;
        test_data[1543] = 33'd5691633262;
        test_addr[1544] = 461;
        test_data[1544] = 33'd583606136;
        test_addr[1545] = 462;
        test_data[1545] = 33'd3772793346;
        test_addr[1546] = 463;
        test_data[1546] = 33'd1274767714;
        test_addr[1547] = 464;
        test_data[1547] = 33'd1701612275;
        test_addr[1548] = 465;
        test_data[1548] = 33'd7435375248;
        test_addr[1549] = 466;
        test_data[1549] = 33'd2807963646;
        test_addr[1550] = 467;
        test_data[1550] = 33'd962725890;
        test_addr[1551] = 468;
        test_data[1551] = 33'd2873278775;
        test_addr[1552] = 469;
        test_data[1552] = 33'd8403157223;
        test_addr[1553] = 470;
        test_data[1553] = 33'd1183712898;
        test_addr[1554] = 471;
        test_data[1554] = 33'd5340606591;
        test_addr[1555] = 472;
        test_data[1555] = 33'd5668775496;
        test_addr[1556] = 473;
        test_data[1556] = 33'd2376303146;
        test_addr[1557] = 474;
        test_data[1557] = 33'd7540287353;
        test_addr[1558] = 694;
        test_data[1558] = 33'd7359557132;
        test_addr[1559] = 695;
        test_data[1559] = 33'd2233471613;
        test_addr[1560] = 696;
        test_data[1560] = 33'd510585055;
        test_addr[1561] = 697;
        test_data[1561] = 33'd241466137;
        test_addr[1562] = 698;
        test_data[1562] = 33'd1941058159;
        test_addr[1563] = 643;
        test_data[1563] = 33'd3900038649;
        test_addr[1564] = 699;
        test_data[1564] = 33'd7198726069;
        test_addr[1565] = 700;
        test_data[1565] = 33'd4290278596;
        test_addr[1566] = 701;
        test_data[1566] = 33'd4872797988;
        test_addr[1567] = 702;
        test_data[1567] = 33'd1769260887;
        test_addr[1568] = 703;
        test_data[1568] = 33'd892604545;
        test_addr[1569] = 704;
        test_data[1569] = 33'd8264563783;
        test_addr[1570] = 705;
        test_data[1570] = 33'd2046342139;
        test_addr[1571] = 706;
        test_data[1571] = 33'd1271505191;
        test_addr[1572] = 707;
        test_data[1572] = 33'd986566342;
        test_addr[1573] = 708;
        test_data[1573] = 33'd2576467063;
        test_addr[1574] = 364;
        test_data[1574] = 33'd4047546126;
        test_addr[1575] = 365;
        test_data[1575] = 33'd1008210114;
        test_addr[1576] = 366;
        test_data[1576] = 33'd2115114658;
        test_addr[1577] = 367;
        test_data[1577] = 33'd916394114;
        test_addr[1578] = 368;
        test_data[1578] = 33'd1550869304;
        test_addr[1579] = 369;
        test_data[1579] = 33'd2180183636;
        test_addr[1580] = 370;
        test_data[1580] = 33'd8334036800;
        test_addr[1581] = 371;
        test_data[1581] = 33'd1796770481;
        test_addr[1582] = 372;
        test_data[1582] = 33'd7895670969;
        test_addr[1583] = 709;
        test_data[1583] = 33'd83794451;
        test_addr[1584] = 710;
        test_data[1584] = 33'd7510558045;
        test_addr[1585] = 711;
        test_data[1585] = 33'd3928838089;
        test_addr[1586] = 712;
        test_data[1586] = 33'd6550220011;
        test_addr[1587] = 713;
        test_data[1587] = 33'd3261845956;
        test_addr[1588] = 714;
        test_data[1588] = 33'd4226705526;
        test_addr[1589] = 715;
        test_data[1589] = 33'd3264214500;
        test_addr[1590] = 833;
        test_data[1590] = 33'd4739310282;
        test_addr[1591] = 834;
        test_data[1591] = 33'd7415941274;
        test_addr[1592] = 835;
        test_data[1592] = 33'd461723609;
        test_addr[1593] = 836;
        test_data[1593] = 33'd433352462;
        test_addr[1594] = 716;
        test_data[1594] = 33'd5122416793;
        test_addr[1595] = 515;
        test_data[1595] = 33'd4175963926;
        test_addr[1596] = 717;
        test_data[1596] = 33'd3532130073;
        test_addr[1597] = 718;
        test_data[1597] = 33'd2494614555;
        test_addr[1598] = 719;
        test_data[1598] = 33'd6619450958;
        test_addr[1599] = 720;
        test_data[1599] = 33'd2104937406;
        test_addr[1600] = 721;
        test_data[1600] = 33'd5423720668;
        test_addr[1601] = 722;
        test_data[1601] = 33'd2657954045;
        test_addr[1602] = 723;
        test_data[1602] = 33'd3748128516;
        test_addr[1603] = 724;
        test_data[1603] = 33'd3564607404;
        test_addr[1604] = 725;
        test_data[1604] = 33'd5953913519;
        test_addr[1605] = 726;
        test_data[1605] = 33'd6604316082;
        test_addr[1606] = 727;
        test_data[1606] = 33'd7766647245;
        test_addr[1607] = 728;
        test_data[1607] = 33'd1284317235;
        test_addr[1608] = 729;
        test_data[1608] = 33'd919345546;
        test_addr[1609] = 730;
        test_data[1609] = 33'd4067928788;
        test_addr[1610] = 731;
        test_data[1610] = 33'd1353510671;
        test_addr[1611] = 732;
        test_data[1611] = 33'd3538750273;
        test_addr[1612] = 733;
        test_data[1612] = 33'd4934107819;
        test_addr[1613] = 734;
        test_data[1613] = 33'd6938553628;
        test_addr[1614] = 735;
        test_data[1614] = 33'd8371444322;
        test_addr[1615] = 736;
        test_data[1615] = 33'd7014823001;
        test_addr[1616] = 737;
        test_data[1616] = 33'd3370945044;
        test_addr[1617] = 738;
        test_data[1617] = 33'd4794622059;
        test_addr[1618] = 739;
        test_data[1618] = 33'd3426545964;
        test_addr[1619] = 740;
        test_data[1619] = 33'd3233147737;
        test_addr[1620] = 741;
        test_data[1620] = 33'd1810153704;
        test_addr[1621] = 742;
        test_data[1621] = 33'd2878401245;
        test_addr[1622] = 545;
        test_data[1622] = 33'd1629998795;
        test_addr[1623] = 546;
        test_data[1623] = 33'd3814328262;
        test_addr[1624] = 547;
        test_data[1624] = 33'd5804834311;
        test_addr[1625] = 548;
        test_data[1625] = 33'd1180199925;
        test_addr[1626] = 549;
        test_data[1626] = 33'd2477350668;
        test_addr[1627] = 550;
        test_data[1627] = 33'd4589490729;
        test_addr[1628] = 551;
        test_data[1628] = 33'd318746959;
        test_addr[1629] = 552;
        test_data[1629] = 33'd2228775572;
        test_addr[1630] = 553;
        test_data[1630] = 33'd6539835559;
        test_addr[1631] = 554;
        test_data[1631] = 33'd3262924390;
        test_addr[1632] = 555;
        test_data[1632] = 33'd449821878;
        test_addr[1633] = 743;
        test_data[1633] = 33'd5206577861;
        test_addr[1634] = 744;
        test_data[1634] = 33'd3214813081;
        test_addr[1635] = 745;
        test_data[1635] = 33'd7599700964;
        test_addr[1636] = 746;
        test_data[1636] = 33'd5570670412;
        test_addr[1637] = 747;
        test_data[1637] = 33'd2220256742;
        test_addr[1638] = 748;
        test_data[1638] = 33'd1521829790;
        test_addr[1639] = 749;
        test_data[1639] = 33'd3952188244;
        test_addr[1640] = 750;
        test_data[1640] = 33'd7894335115;
        test_addr[1641] = 751;
        test_data[1641] = 33'd3419461017;
        test_addr[1642] = 752;
        test_data[1642] = 33'd467983000;
        test_addr[1643] = 753;
        test_data[1643] = 33'd4101479975;
        test_addr[1644] = 754;
        test_data[1644] = 33'd2930249500;
        test_addr[1645] = 755;
        test_data[1645] = 33'd227107951;
        test_addr[1646] = 756;
        test_data[1646] = 33'd1338030971;
        test_addr[1647] = 757;
        test_data[1647] = 33'd2619751839;
        test_addr[1648] = 758;
        test_data[1648] = 33'd4562143389;
        test_addr[1649] = 759;
        test_data[1649] = 33'd1446998705;
        test_addr[1650] = 760;
        test_data[1650] = 33'd3811051108;
        test_addr[1651] = 761;
        test_data[1651] = 33'd5989830610;
        test_addr[1652] = 762;
        test_data[1652] = 33'd3993692466;
        test_addr[1653] = 763;
        test_data[1653] = 33'd930239523;
        test_addr[1654] = 764;
        test_data[1654] = 33'd6603898777;
        test_addr[1655] = 765;
        test_data[1655] = 33'd8502460255;
        test_addr[1656] = 766;
        test_data[1656] = 33'd910969802;
        test_addr[1657] = 767;
        test_data[1657] = 33'd2089824228;
        test_addr[1658] = 768;
        test_data[1658] = 33'd4646774037;
        test_addr[1659] = 769;
        test_data[1659] = 33'd3880414256;
        test_addr[1660] = 770;
        test_data[1660] = 33'd317508578;
        test_addr[1661] = 771;
        test_data[1661] = 33'd7930569419;
        test_addr[1662] = 772;
        test_data[1662] = 33'd1620593328;
        test_addr[1663] = 773;
        test_data[1663] = 33'd256807720;
        test_addr[1664] = 774;
        test_data[1664] = 33'd9534195;
        test_addr[1665] = 775;
        test_data[1665] = 33'd5324830943;
        test_addr[1666] = 776;
        test_data[1666] = 33'd3596983855;
        test_addr[1667] = 647;
        test_data[1667] = 33'd4792275722;
        test_addr[1668] = 648;
        test_data[1668] = 33'd7121756174;
        test_addr[1669] = 649;
        test_data[1669] = 33'd4680511418;
        test_addr[1670] = 777;
        test_data[1670] = 33'd3617657151;
        test_addr[1671] = 778;
        test_data[1671] = 33'd1257411684;
        test_addr[1672] = 571;
        test_data[1672] = 33'd4869237358;
        test_addr[1673] = 572;
        test_data[1673] = 33'd2320974549;
        test_addr[1674] = 573;
        test_data[1674] = 33'd5242795131;
        test_addr[1675] = 779;
        test_data[1675] = 33'd6427914744;
        test_addr[1676] = 634;
        test_data[1676] = 33'd954992338;
        test_addr[1677] = 635;
        test_data[1677] = 33'd3974692757;
        test_addr[1678] = 636;
        test_data[1678] = 33'd4218479966;
        test_addr[1679] = 637;
        test_data[1679] = 33'd3795165725;
        test_addr[1680] = 638;
        test_data[1680] = 33'd881995127;
        test_addr[1681] = 639;
        test_data[1681] = 33'd2250332921;
        test_addr[1682] = 640;
        test_data[1682] = 33'd561070447;
        test_addr[1683] = 641;
        test_data[1683] = 33'd2087204287;
        test_addr[1684] = 642;
        test_data[1684] = 33'd771630044;
        test_addr[1685] = 643;
        test_data[1685] = 33'd3900038649;
        test_addr[1686] = 644;
        test_data[1686] = 33'd3175733827;
        test_addr[1687] = 645;
        test_data[1687] = 33'd4069788299;
        test_addr[1688] = 780;
        test_data[1688] = 33'd1167957788;
        test_addr[1689] = 781;
        test_data[1689] = 33'd1128514710;
        test_addr[1690] = 782;
        test_data[1690] = 33'd2652390457;
        test_addr[1691] = 783;
        test_data[1691] = 33'd5776899834;
        test_addr[1692] = 784;
        test_data[1692] = 33'd3365509421;
        test_addr[1693] = 785;
        test_data[1693] = 33'd4360038821;
        test_addr[1694] = 786;
        test_data[1694] = 33'd3695516988;
        test_addr[1695] = 787;
        test_data[1695] = 33'd828291663;
        test_addr[1696] = 788;
        test_data[1696] = 33'd1105670773;
        test_addr[1697] = 789;
        test_data[1697] = 33'd911008138;
        test_addr[1698] = 790;
        test_data[1698] = 33'd1470099950;
        test_addr[1699] = 791;
        test_data[1699] = 33'd5892966168;
        test_addr[1700] = 792;
        test_data[1700] = 33'd5089624170;
        test_addr[1701] = 793;
        test_data[1701] = 33'd1321282978;
        test_addr[1702] = 794;
        test_data[1702] = 33'd5729956780;
        test_addr[1703] = 795;
        test_data[1703] = 33'd5865181433;
        test_addr[1704] = 796;
        test_data[1704] = 33'd2646907564;
        test_addr[1705] = 797;
        test_data[1705] = 33'd99933581;
        test_addr[1706] = 134;
        test_data[1706] = 33'd7281480161;
        test_addr[1707] = 135;
        test_data[1707] = 33'd1960021159;
        test_addr[1708] = 136;
        test_data[1708] = 33'd3552771192;
        test_addr[1709] = 137;
        test_data[1709] = 33'd8325876202;
        test_addr[1710] = 138;
        test_data[1710] = 33'd6412243605;
        test_addr[1711] = 798;
        test_data[1711] = 33'd3837150160;
        test_addr[1712] = 799;
        test_data[1712] = 33'd3441245320;
        test_addr[1713] = 800;
        test_data[1713] = 33'd6952853902;
        test_addr[1714] = 801;
        test_data[1714] = 33'd1686375627;
        test_addr[1715] = 802;
        test_data[1715] = 33'd4239473607;
        test_addr[1716] = 803;
        test_data[1716] = 33'd7634248285;
        test_addr[1717] = 804;
        test_data[1717] = 33'd1315671584;
        test_addr[1718] = 805;
        test_data[1718] = 33'd3455870968;
        test_addr[1719] = 806;
        test_data[1719] = 33'd1359101487;
        test_addr[1720] = 807;
        test_data[1720] = 33'd540490609;
        test_addr[1721] = 808;
        test_data[1721] = 33'd4179863201;
        test_addr[1722] = 809;
        test_data[1722] = 33'd8061903279;
        test_addr[1723] = 810;
        test_data[1723] = 33'd8350996439;
        test_addr[1724] = 225;
        test_data[1724] = 33'd206097148;
        test_addr[1725] = 226;
        test_data[1725] = 33'd2883781805;
        test_addr[1726] = 227;
        test_data[1726] = 33'd355985290;
        test_addr[1727] = 228;
        test_data[1727] = 33'd4334309053;
        test_addr[1728] = 229;
        test_data[1728] = 33'd845232644;
        test_addr[1729] = 230;
        test_data[1729] = 33'd4730375106;
        test_addr[1730] = 231;
        test_data[1730] = 33'd164270080;
        test_addr[1731] = 232;
        test_data[1731] = 33'd111204031;
        test_addr[1732] = 233;
        test_data[1732] = 33'd2304627638;
        test_addr[1733] = 234;
        test_data[1733] = 33'd7006710871;
        test_addr[1734] = 235;
        test_data[1734] = 33'd1995153683;
        test_addr[1735] = 236;
        test_data[1735] = 33'd3308823479;
        test_addr[1736] = 237;
        test_data[1736] = 33'd5990711261;
        test_addr[1737] = 238;
        test_data[1737] = 33'd6325111245;
        test_addr[1738] = 811;
        test_data[1738] = 33'd4552623601;
        test_addr[1739] = 812;
        test_data[1739] = 33'd3444397451;
        test_addr[1740] = 813;
        test_data[1740] = 33'd3209556232;
        test_addr[1741] = 814;
        test_data[1741] = 33'd3061961020;
        test_addr[1742] = 815;
        test_data[1742] = 33'd99083937;
        test_addr[1743] = 816;
        test_data[1743] = 33'd3371550778;
        test_addr[1744] = 817;
        test_data[1744] = 33'd7521436164;
        test_addr[1745] = 818;
        test_data[1745] = 33'd4841791642;
        test_addr[1746] = 819;
        test_data[1746] = 33'd7949724091;
        test_addr[1747] = 820;
        test_data[1747] = 33'd1650346404;
        test_addr[1748] = 821;
        test_data[1748] = 33'd971615072;
        test_addr[1749] = 822;
        test_data[1749] = 33'd7116640242;
        test_addr[1750] = 823;
        test_data[1750] = 33'd532265002;
        test_addr[1751] = 397;
        test_data[1751] = 33'd3874668741;
        test_addr[1752] = 398;
        test_data[1752] = 33'd2124586123;
        test_addr[1753] = 399;
        test_data[1753] = 33'd7367503479;
        test_addr[1754] = 400;
        test_data[1754] = 33'd6555915342;
        test_addr[1755] = 401;
        test_data[1755] = 33'd5272491017;
        test_addr[1756] = 402;
        test_data[1756] = 33'd246986956;
        test_addr[1757] = 403;
        test_data[1757] = 33'd603897780;
        test_addr[1758] = 404;
        test_data[1758] = 33'd284306586;
        test_addr[1759] = 405;
        test_data[1759] = 33'd7476641818;
        test_addr[1760] = 406;
        test_data[1760] = 33'd2830641639;
        test_addr[1761] = 407;
        test_data[1761] = 33'd7604336461;
        test_addr[1762] = 408;
        test_data[1762] = 33'd7827813012;
        test_addr[1763] = 409;
        test_data[1763] = 33'd6003201581;
        test_addr[1764] = 410;
        test_data[1764] = 33'd3422075366;
        test_addr[1765] = 411;
        test_data[1765] = 33'd3626126882;
        test_addr[1766] = 412;
        test_data[1766] = 33'd5801849477;
        test_addr[1767] = 413;
        test_data[1767] = 33'd2482816989;
        test_addr[1768] = 824;
        test_data[1768] = 33'd3204893334;
        test_addr[1769] = 825;
        test_data[1769] = 33'd7535788355;
        test_addr[1770] = 826;
        test_data[1770] = 33'd2805664193;
        test_addr[1771] = 827;
        test_data[1771] = 33'd1406447338;
        test_addr[1772] = 828;
        test_data[1772] = 33'd1271401654;
        test_addr[1773] = 829;
        test_data[1773] = 33'd7220600844;
        test_addr[1774] = 830;
        test_data[1774] = 33'd8483735687;
        test_addr[1775] = 831;
        test_data[1775] = 33'd4718344998;
        test_addr[1776] = 832;
        test_data[1776] = 33'd6046332013;
        test_addr[1777] = 833;
        test_data[1777] = 33'd444342986;
        test_addr[1778] = 834;
        test_data[1778] = 33'd3120973978;
        test_addr[1779] = 835;
        test_data[1779] = 33'd461723609;
        test_addr[1780] = 836;
        test_data[1780] = 33'd433352462;
        test_addr[1781] = 837;
        test_data[1781] = 33'd1959645325;
        test_addr[1782] = 838;
        test_data[1782] = 33'd3573850885;
        test_addr[1783] = 839;
        test_data[1783] = 33'd1323733114;
        test_addr[1784] = 577;
        test_data[1784] = 33'd1793952775;
        test_addr[1785] = 578;
        test_data[1785] = 33'd3196294421;
        test_addr[1786] = 579;
        test_data[1786] = 33'd1094013198;
        test_addr[1787] = 580;
        test_data[1787] = 33'd1233267658;
        test_addr[1788] = 581;
        test_data[1788] = 33'd4657789767;
        test_addr[1789] = 582;
        test_data[1789] = 33'd3179541911;
        test_addr[1790] = 583;
        test_data[1790] = 33'd2231704842;
        test_addr[1791] = 584;
        test_data[1791] = 33'd1490217735;
        test_addr[1792] = 585;
        test_data[1792] = 33'd1270660057;
        test_addr[1793] = 586;
        test_data[1793] = 33'd1844798620;
        test_addr[1794] = 587;
        test_data[1794] = 33'd5661226171;
        test_addr[1795] = 588;
        test_data[1795] = 33'd1893529001;
        test_addr[1796] = 589;
        test_data[1796] = 33'd3514985912;
        test_addr[1797] = 590;
        test_data[1797] = 33'd2083229337;
        test_addr[1798] = 591;
        test_data[1798] = 33'd8290171892;
        test_addr[1799] = 592;
        test_data[1799] = 33'd6271769546;
        test_addr[1800] = 593;
        test_data[1800] = 33'd704520665;
        test_addr[1801] = 594;
        test_data[1801] = 33'd499927349;
        test_addr[1802] = 595;
        test_data[1802] = 33'd4658576337;
        test_addr[1803] = 596;
        test_data[1803] = 33'd2164998835;
        test_addr[1804] = 597;
        test_data[1804] = 33'd4269111753;
        test_addr[1805] = 598;
        test_data[1805] = 33'd3698561184;
        test_addr[1806] = 599;
        test_data[1806] = 33'd2621666958;
        test_addr[1807] = 600;
        test_data[1807] = 33'd1029049725;
        test_addr[1808] = 601;
        test_data[1808] = 33'd647592843;
        test_addr[1809] = 602;
        test_data[1809] = 33'd4563852132;
        test_addr[1810] = 603;
        test_data[1810] = 33'd3565486424;
        test_addr[1811] = 604;
        test_data[1811] = 33'd7443273777;
        test_addr[1812] = 605;
        test_data[1812] = 33'd4068052147;
        test_addr[1813] = 606;
        test_data[1813] = 33'd906696308;
        test_addr[1814] = 607;
        test_data[1814] = 33'd5620450195;
        test_addr[1815] = 608;
        test_data[1815] = 33'd3635138265;
        test_addr[1816] = 609;
        test_data[1816] = 33'd2142050983;
        test_addr[1817] = 840;
        test_data[1817] = 33'd462945108;
        test_addr[1818] = 841;
        test_data[1818] = 33'd729735648;
        test_addr[1819] = 842;
        test_data[1819] = 33'd3905935845;
        test_addr[1820] = 843;
        test_data[1820] = 33'd64812169;
        test_addr[1821] = 844;
        test_data[1821] = 33'd1905889562;
        test_addr[1822] = 845;
        test_data[1822] = 33'd4716021179;
        test_addr[1823] = 846;
        test_data[1823] = 33'd3157279990;
        test_addr[1824] = 847;
        test_data[1824] = 33'd4178636307;
        test_addr[1825] = 848;
        test_data[1825] = 33'd1091101872;
        test_addr[1826] = 849;
        test_data[1826] = 33'd2875037109;
        test_addr[1827] = 850;
        test_data[1827] = 33'd1086596891;
        test_addr[1828] = 851;
        test_data[1828] = 33'd30109657;
        test_addr[1829] = 852;
        test_data[1829] = 33'd6824448436;
        test_addr[1830] = 853;
        test_data[1830] = 33'd5848566463;
        test_addr[1831] = 854;
        test_data[1831] = 33'd6562141206;
        test_addr[1832] = 855;
        test_data[1832] = 33'd3155227187;
        test_addr[1833] = 856;
        test_data[1833] = 33'd2735570664;
        test_addr[1834] = 857;
        test_data[1834] = 33'd5978025865;
        test_addr[1835] = 858;
        test_data[1835] = 33'd3668307118;
        test_addr[1836] = 859;
        test_data[1836] = 33'd790427723;
        test_addr[1837] = 860;
        test_data[1837] = 33'd2040878775;
        test_addr[1838] = 861;
        test_data[1838] = 33'd2853075293;
        test_addr[1839] = 862;
        test_data[1839] = 33'd3234096972;
        test_addr[1840] = 339;
        test_data[1840] = 33'd4509445827;
        test_addr[1841] = 340;
        test_data[1841] = 33'd451413948;
        test_addr[1842] = 341;
        test_data[1842] = 33'd5037414763;
        test_addr[1843] = 342;
        test_data[1843] = 33'd5921216805;
        test_addr[1844] = 343;
        test_data[1844] = 33'd5693607392;
        test_addr[1845] = 344;
        test_data[1845] = 33'd281373290;
        test_addr[1846] = 863;
        test_data[1846] = 33'd983979571;
        test_addr[1847] = 864;
        test_data[1847] = 33'd2537001022;
        test_addr[1848] = 513;
        test_data[1848] = 33'd3832833658;
        test_addr[1849] = 514;
        test_data[1849] = 33'd1741233038;
        test_addr[1850] = 865;
        test_data[1850] = 33'd7304379496;
        test_addr[1851] = 866;
        test_data[1851] = 33'd2528451676;
        test_addr[1852] = 187;
        test_data[1852] = 33'd8572842172;
        test_addr[1853] = 867;
        test_data[1853] = 33'd4195620311;
        test_addr[1854] = 868;
        test_data[1854] = 33'd749785393;
        test_addr[1855] = 869;
        test_data[1855] = 33'd3921532732;
        test_addr[1856] = 870;
        test_data[1856] = 33'd7440125811;
        test_addr[1857] = 871;
        test_data[1857] = 33'd3229558777;
        test_addr[1858] = 872;
        test_data[1858] = 33'd4656759110;
        test_addr[1859] = 873;
        test_data[1859] = 33'd1520019581;
        test_addr[1860] = 874;
        test_data[1860] = 33'd4813375875;
        test_addr[1861] = 875;
        test_data[1861] = 33'd1778218794;
        test_addr[1862] = 876;
        test_data[1862] = 33'd3812382912;
        test_addr[1863] = 641;
        test_data[1863] = 33'd2087204287;
        test_addr[1864] = 642;
        test_data[1864] = 33'd771630044;
        test_addr[1865] = 643;
        test_data[1865] = 33'd3900038649;
        test_addr[1866] = 644;
        test_data[1866] = 33'd3175733827;
        test_addr[1867] = 877;
        test_data[1867] = 33'd2926156055;
        test_addr[1868] = 878;
        test_data[1868] = 33'd8020475481;
        test_addr[1869] = 879;
        test_data[1869] = 33'd4619439445;
        test_addr[1870] = 880;
        test_data[1870] = 33'd7559541088;
        test_addr[1871] = 881;
        test_data[1871] = 33'd4451175104;
        test_addr[1872] = 535;
        test_data[1872] = 33'd2501250615;
        test_addr[1873] = 536;
        test_data[1873] = 33'd6312695888;
        test_addr[1874] = 537;
        test_data[1874] = 33'd7991570926;
        test_addr[1875] = 538;
        test_data[1875] = 33'd7009801064;
        test_addr[1876] = 539;
        test_data[1876] = 33'd2749828337;
        test_addr[1877] = 540;
        test_data[1877] = 33'd30470061;
        test_addr[1878] = 541;
        test_data[1878] = 33'd2310349212;
        test_addr[1879] = 542;
        test_data[1879] = 33'd2967622748;
        test_addr[1880] = 543;
        test_data[1880] = 33'd298678754;
        test_addr[1881] = 544;
        test_data[1881] = 33'd7250787811;
        test_addr[1882] = 545;
        test_data[1882] = 33'd1629998795;
        test_addr[1883] = 546;
        test_data[1883] = 33'd5579341168;
        test_addr[1884] = 547;
        test_data[1884] = 33'd6433181043;
        test_addr[1885] = 548;
        test_data[1885] = 33'd8575742989;
        test_addr[1886] = 882;
        test_data[1886] = 33'd7864792130;
        test_addr[1887] = 883;
        test_data[1887] = 33'd4733896684;
        test_addr[1888] = 83;
        test_data[1888] = 33'd176121797;
        test_addr[1889] = 84;
        test_data[1889] = 33'd389769389;
        test_addr[1890] = 85;
        test_data[1890] = 33'd3382751907;
        test_addr[1891] = 884;
        test_data[1891] = 33'd700616692;
        test_addr[1892] = 885;
        test_data[1892] = 33'd3458389258;
        test_addr[1893] = 886;
        test_data[1893] = 33'd7113117625;
        test_addr[1894] = 887;
        test_data[1894] = 33'd2507313658;
        test_addr[1895] = 888;
        test_data[1895] = 33'd397640837;
        test_addr[1896] = 889;
        test_data[1896] = 33'd1528309135;
        test_addr[1897] = 890;
        test_data[1897] = 33'd42358296;
        test_addr[1898] = 175;
        test_data[1898] = 33'd3567745488;
        test_addr[1899] = 891;
        test_data[1899] = 33'd6910032508;
        test_addr[1900] = 892;
        test_data[1900] = 33'd5080764799;
        test_addr[1901] = 893;
        test_data[1901] = 33'd4472798289;
        test_addr[1902] = 811;
        test_data[1902] = 33'd257656305;
        test_addr[1903] = 812;
        test_data[1903] = 33'd4793032381;
        test_addr[1904] = 813;
        test_data[1904] = 33'd3209556232;
        test_addr[1905] = 814;
        test_data[1905] = 33'd8299652681;
        test_addr[1906] = 815;
        test_data[1906] = 33'd4405663113;
        test_addr[1907] = 816;
        test_data[1907] = 33'd4768992363;
        test_addr[1908] = 817;
        test_data[1908] = 33'd5181838644;
        test_addr[1909] = 818;
        test_data[1909] = 33'd546824346;
        test_addr[1910] = 819;
        test_data[1910] = 33'd5465227510;
        test_addr[1911] = 820;
        test_data[1911] = 33'd1650346404;
        test_addr[1912] = 821;
        test_data[1912] = 33'd971615072;
        test_addr[1913] = 822;
        test_data[1913] = 33'd2821672946;
        test_addr[1914] = 823;
        test_data[1914] = 33'd532265002;
        test_addr[1915] = 824;
        test_data[1915] = 33'd3204893334;
        test_addr[1916] = 825;
        test_data[1916] = 33'd3240821059;
        test_addr[1917] = 826;
        test_data[1917] = 33'd7931402239;
        test_addr[1918] = 827;
        test_data[1918] = 33'd1406447338;
        test_addr[1919] = 828;
        test_data[1919] = 33'd1271401654;
        test_addr[1920] = 829;
        test_data[1920] = 33'd4682295617;
        test_addr[1921] = 830;
        test_data[1921] = 33'd4188768391;
        test_addr[1922] = 831;
        test_data[1922] = 33'd423377702;
        test_addr[1923] = 832;
        test_data[1923] = 33'd8233945145;
        test_addr[1924] = 833;
        test_data[1924] = 33'd444342986;
        test_addr[1925] = 834;
        test_data[1925] = 33'd7628206370;
        test_addr[1926] = 835;
        test_data[1926] = 33'd461723609;
        test_addr[1927] = 836;
        test_data[1927] = 33'd433352462;
        test_addr[1928] = 837;
        test_data[1928] = 33'd1959645325;
        test_addr[1929] = 838;
        test_data[1929] = 33'd3573850885;
        test_addr[1930] = 839;
        test_data[1930] = 33'd1323733114;
        test_addr[1931] = 894;
        test_data[1931] = 33'd585438621;
        test_addr[1932] = 895;
        test_data[1932] = 33'd3072952231;
        test_addr[1933] = 896;
        test_data[1933] = 33'd819431204;
        test_addr[1934] = 897;
        test_data[1934] = 33'd268761716;
        test_addr[1935] = 898;
        test_data[1935] = 33'd1775297931;
        test_addr[1936] = 899;
        test_data[1936] = 33'd8513902736;
        test_addr[1937] = 900;
        test_data[1937] = 33'd2081706384;
        test_addr[1938] = 220;
        test_data[1938] = 33'd728361109;
        test_addr[1939] = 221;
        test_data[1939] = 33'd1780024880;
        test_addr[1940] = 222;
        test_data[1940] = 33'd4233733742;
        test_addr[1941] = 223;
        test_data[1941] = 33'd3770350222;
        test_addr[1942] = 224;
        test_data[1942] = 33'd3332430587;
        test_addr[1943] = 225;
        test_data[1943] = 33'd206097148;
        test_addr[1944] = 901;
        test_data[1944] = 33'd1604865859;
        test_addr[1945] = 902;
        test_data[1945] = 33'd8057080010;
        test_addr[1946] = 903;
        test_data[1946] = 33'd486481265;
        test_addr[1947] = 904;
        test_data[1947] = 33'd299855562;
        test_addr[1948] = 905;
        test_data[1948] = 33'd1328078859;
        test_addr[1949] = 906;
        test_data[1949] = 33'd8302344222;
        test_addr[1950] = 907;
        test_data[1950] = 33'd1829404985;
        test_addr[1951] = 908;
        test_data[1951] = 33'd3676688916;
        test_addr[1952] = 909;
        test_data[1952] = 33'd6886092515;
        test_addr[1953] = 910;
        test_data[1953] = 33'd6689410811;
        test_addr[1954] = 911;
        test_data[1954] = 33'd806648968;
        test_addr[1955] = 912;
        test_data[1955] = 33'd5311297690;
        test_addr[1956] = 913;
        test_data[1956] = 33'd858191111;
        test_addr[1957] = 1018;
        test_data[1957] = 33'd2750972131;
        test_addr[1958] = 1019;
        test_data[1958] = 33'd6356435954;
        test_addr[1959] = 1020;
        test_data[1959] = 33'd6514373451;
        test_addr[1960] = 1021;
        test_data[1960] = 33'd7300244544;
        test_addr[1961] = 1022;
        test_data[1961] = 33'd2746665182;
        test_addr[1962] = 1023;
        test_data[1962] = 33'd4086440552;
        test_addr[1963] = 0;
        test_data[1963] = 33'd1870585436;
        test_addr[1964] = 914;
        test_data[1964] = 33'd4191420171;
        test_addr[1965] = 915;
        test_data[1965] = 33'd8054869188;
        test_addr[1966] = 916;
        test_data[1966] = 33'd936149391;
        test_addr[1967] = 917;
        test_data[1967] = 33'd7819878378;
        test_addr[1968] = 945;
        test_data[1968] = 33'd5637592309;
        test_addr[1969] = 946;
        test_data[1969] = 33'd1984305920;
        test_addr[1970] = 918;
        test_data[1970] = 33'd3381071146;
        test_addr[1971] = 919;
        test_data[1971] = 33'd632463510;
        test_addr[1972] = 920;
        test_data[1972] = 33'd7929007260;
        test_addr[1973] = 921;
        test_data[1973] = 33'd7287081892;
        test_addr[1974] = 922;
        test_data[1974] = 33'd2267903388;
        test_addr[1975] = 923;
        test_data[1975] = 33'd3334114139;
        test_addr[1976] = 979;
        test_data[1976] = 33'd3552257411;
        test_addr[1977] = 980;
        test_data[1977] = 33'd3721886817;
        test_addr[1978] = 981;
        test_data[1978] = 33'd166781239;
        test_addr[1979] = 982;
        test_data[1979] = 33'd2064422908;
        test_addr[1980] = 924;
        test_data[1980] = 33'd2084629605;
        test_addr[1981] = 925;
        test_data[1981] = 33'd2610089944;
        test_addr[1982] = 926;
        test_data[1982] = 33'd7440282351;
        test_addr[1983] = 927;
        test_data[1983] = 33'd425505923;
        test_addr[1984] = 928;
        test_data[1984] = 33'd1778724627;
        test_addr[1985] = 929;
        test_data[1985] = 33'd8060946427;
        test_addr[1986] = 930;
        test_data[1986] = 33'd1564872363;
        test_addr[1987] = 931;
        test_data[1987] = 33'd4191689811;
        test_addr[1988] = 932;
        test_data[1988] = 33'd7973407690;
        test_addr[1989] = 300;
        test_data[1989] = 33'd6174988878;
        test_addr[1990] = 301;
        test_data[1990] = 33'd779647779;
        test_addr[1991] = 302;
        test_data[1991] = 33'd2759854552;
        test_addr[1992] = 303;
        test_data[1992] = 33'd4351636344;
        test_addr[1993] = 304;
        test_data[1993] = 33'd4755795012;
        test_addr[1994] = 305;
        test_data[1994] = 33'd1866235150;
        test_addr[1995] = 306;
        test_data[1995] = 33'd1400119106;
        test_addr[1996] = 307;
        test_data[1996] = 33'd4593616462;
        test_addr[1997] = 308;
        test_data[1997] = 33'd2611705428;
        test_addr[1998] = 309;
        test_data[1998] = 33'd3941608837;
        test_addr[1999] = 310;
        test_data[1999] = 33'd3094631771;
        test_addr[2000] = 311;
        test_data[2000] = 33'd1449524691;
        test_addr[2001] = 312;
        test_data[2001] = 33'd240548675;
        test_addr[2002] = 313;
        test_data[2002] = 33'd3069166694;
        test_addr[2003] = 314;
        test_data[2003] = 33'd2141065806;
        test_addr[2004] = 315;
        test_data[2004] = 33'd3309303920;
        test_addr[2005] = 933;
        test_data[2005] = 33'd170108847;
        test_addr[2006] = 665;
        test_data[2006] = 33'd6206541747;
        test_addr[2007] = 666;
        test_data[2007] = 33'd8289936758;
        test_addr[2008] = 667;
        test_data[2008] = 33'd3634324503;
        test_addr[2009] = 668;
        test_data[2009] = 33'd6643889209;
        test_addr[2010] = 669;
        test_data[2010] = 33'd100741952;
        test_addr[2011] = 670;
        test_data[2011] = 33'd3197879796;
        test_addr[2012] = 671;
        test_data[2012] = 33'd3754236325;
        test_addr[2013] = 672;
        test_data[2013] = 33'd1411628437;
        test_addr[2014] = 673;
        test_data[2014] = 33'd7786648293;
        test_addr[2015] = 934;
        test_data[2015] = 33'd5624971451;
        test_addr[2016] = 935;
        test_data[2016] = 33'd6268741827;
        test_addr[2017] = 936;
        test_data[2017] = 33'd607348316;
        test_addr[2018] = 937;
        test_data[2018] = 33'd625389764;
        test_addr[2019] = 938;
        test_data[2019] = 33'd4416210223;
        test_addr[2020] = 939;
        test_data[2020] = 33'd349632060;
        test_addr[2021] = 940;
        test_data[2021] = 33'd3211187226;
        test_addr[2022] = 941;
        test_data[2022] = 33'd1460688612;
        test_addr[2023] = 942;
        test_data[2023] = 33'd3185997769;
        test_addr[2024] = 943;
        test_data[2024] = 33'd1653503808;
        test_addr[2025] = 944;
        test_data[2025] = 33'd1934668787;
        test_addr[2026] = 945;
        test_data[2026] = 33'd1342625013;
        test_addr[2027] = 946;
        test_data[2027] = 33'd1984305920;
        test_addr[2028] = 947;
        test_data[2028] = 33'd3397671939;
        test_addr[2029] = 948;
        test_data[2029] = 33'd689974145;
        test_addr[2030] = 949;
        test_data[2030] = 33'd1182899197;
        test_addr[2031] = 950;
        test_data[2031] = 33'd5960325939;
        test_addr[2032] = 951;
        test_data[2032] = 33'd3631193825;
        test_addr[2033] = 952;
        test_data[2033] = 33'd1791314849;
        test_addr[2034] = 953;
        test_data[2034] = 33'd2693867941;
        test_addr[2035] = 954;
        test_data[2035] = 33'd2796648127;
        test_addr[2036] = 955;
        test_data[2036] = 33'd905894982;
        test_addr[2037] = 956;
        test_data[2037] = 33'd90020364;
        test_addr[2038] = 957;
        test_data[2038] = 33'd2991872276;
        test_addr[2039] = 958;
        test_data[2039] = 33'd3447221745;
        test_addr[2040] = 339;
        test_data[2040] = 33'd214478531;
        test_addr[2041] = 340;
        test_data[2041] = 33'd451413948;
        test_addr[2042] = 341;
        test_data[2042] = 33'd742447467;
        test_addr[2043] = 342;
        test_data[2043] = 33'd1626249509;
        test_addr[2044] = 959;
        test_data[2044] = 33'd8089567101;
        test_addr[2045] = 960;
        test_data[2045] = 33'd3497165691;
        test_addr[2046] = 961;
        test_data[2046] = 33'd2075048097;
        test_addr[2047] = 962;
        test_data[2047] = 33'd2765447673;
        test_addr[2048] = 963;
        test_data[2048] = 33'd2156815949;
        test_addr[2049] = 964;
        test_data[2049] = 33'd8230428382;
        test_addr[2050] = 992;
        test_data[2050] = 33'd1625093277;
        test_addr[2051] = 993;
        test_data[2051] = 33'd1150199168;
        test_addr[2052] = 994;
        test_data[2052] = 33'd4788566175;
        test_addr[2053] = 995;
        test_data[2053] = 33'd1594198084;
        test_addr[2054] = 996;
        test_data[2054] = 33'd103670533;
        test_addr[2055] = 997;
        test_data[2055] = 33'd7841847811;
        test_addr[2056] = 998;
        test_data[2056] = 33'd6288932274;
        test_addr[2057] = 965;
        test_data[2057] = 33'd6619240717;
        test_addr[2058] = 960;
        test_data[2058] = 33'd7639929681;
        test_addr[2059] = 961;
        test_data[2059] = 33'd2075048097;
        test_addr[2060] = 962;
        test_data[2060] = 33'd6862146752;
        test_addr[2061] = 963;
        test_data[2061] = 33'd5067628418;
        test_addr[2062] = 964;
        test_data[2062] = 33'd3935461086;
        test_addr[2063] = 966;
        test_data[2063] = 33'd2560894838;
        test_addr[2064] = 967;
        test_data[2064] = 33'd4509235394;
        test_addr[2065] = 968;
        test_data[2065] = 33'd3074093940;
        test_addr[2066] = 969;
        test_data[2066] = 33'd1953469504;
        test_addr[2067] = 970;
        test_data[2067] = 33'd8560430226;
        test_addr[2068] = 971;
        test_data[2068] = 33'd1365898262;
        test_addr[2069] = 972;
        test_data[2069] = 33'd6676586602;
        test_addr[2070] = 973;
        test_data[2070] = 33'd5728811561;
        test_addr[2071] = 974;
        test_data[2071] = 33'd7258037960;
        test_addr[2072] = 975;
        test_data[2072] = 33'd900993035;
        test_addr[2073] = 976;
        test_data[2073] = 33'd888555328;
        test_addr[2074] = 977;
        test_data[2074] = 33'd5662061317;
        test_addr[2075] = 90;
        test_data[2075] = 33'd548807498;
        test_addr[2076] = 91;
        test_data[2076] = 33'd5789302439;
        test_addr[2077] = 92;
        test_data[2077] = 33'd4105109197;
        test_addr[2078] = 93;
        test_data[2078] = 33'd284207449;
        test_addr[2079] = 94;
        test_data[2079] = 33'd8310437457;
        test_addr[2080] = 95;
        test_data[2080] = 33'd767116640;
        test_addr[2081] = 978;
        test_data[2081] = 33'd4907373996;
        test_addr[2082] = 979;
        test_data[2082] = 33'd5342488869;
        test_addr[2083] = 980;
        test_data[2083] = 33'd3721886817;
        test_addr[2084] = 981;
        test_data[2084] = 33'd166781239;
        test_addr[2085] = 96;
        test_data[2085] = 33'd5720597339;
        test_addr[2086] = 97;
        test_data[2086] = 33'd7474211596;
        test_addr[2087] = 98;
        test_data[2087] = 33'd5331022734;
        test_addr[2088] = 99;
        test_data[2088] = 33'd7839220164;
        test_addr[2089] = 100;
        test_data[2089] = 33'd5853096927;
        test_addr[2090] = 101;
        test_data[2090] = 33'd6483585906;
        test_addr[2091] = 102;
        test_data[2091] = 33'd3632082374;
        test_addr[2092] = 103;
        test_data[2092] = 33'd2907570000;
        test_addr[2093] = 104;
        test_data[2093] = 33'd2404063296;
        test_addr[2094] = 105;
        test_data[2094] = 33'd1914703890;
        test_addr[2095] = 106;
        test_data[2095] = 33'd568746040;
        test_addr[2096] = 107;
        test_data[2096] = 33'd2329785644;
        test_addr[2097] = 108;
        test_data[2097] = 33'd3133920479;
        test_addr[2098] = 109;
        test_data[2098] = 33'd2828290416;
        test_addr[2099] = 110;
        test_data[2099] = 33'd8212224405;
        test_addr[2100] = 111;
        test_data[2100] = 33'd7776118917;
        test_addr[2101] = 112;
        test_data[2101] = 33'd1611235687;
        test_addr[2102] = 113;
        test_data[2102] = 33'd8213424307;
        test_addr[2103] = 114;
        test_data[2103] = 33'd6539273879;
        test_addr[2104] = 115;
        test_data[2104] = 33'd1862517686;
        test_addr[2105] = 116;
        test_data[2105] = 33'd1148833960;
        test_addr[2106] = 117;
        test_data[2106] = 33'd6967271051;
        test_addr[2107] = 118;
        test_data[2107] = 33'd4686693002;
        test_addr[2108] = 119;
        test_data[2108] = 33'd2989373656;
        test_addr[2109] = 120;
        test_data[2109] = 33'd7904871636;
        test_addr[2110] = 121;
        test_data[2110] = 33'd371426538;
        test_addr[2111] = 122;
        test_data[2111] = 33'd1367201542;
        test_addr[2112] = 123;
        test_data[2112] = 33'd313859363;
        test_addr[2113] = 124;
        test_data[2113] = 33'd4840436137;
        test_addr[2114] = 982;
        test_data[2114] = 33'd2064422908;
        test_addr[2115] = 983;
        test_data[2115] = 33'd5535518258;
        test_addr[2116] = 984;
        test_data[2116] = 33'd447706912;
        test_addr[2117] = 985;
        test_data[2117] = 33'd6721021472;
        test_addr[2118] = 986;
        test_data[2118] = 33'd8293901458;
        test_addr[2119] = 987;
        test_data[2119] = 33'd6457596556;
        test_addr[2120] = 988;
        test_data[2120] = 33'd1189533474;
        test_addr[2121] = 989;
        test_data[2121] = 33'd1658312967;
        test_addr[2122] = 990;
        test_data[2122] = 33'd431413773;
        test_addr[2123] = 333;
        test_data[2123] = 33'd1462324255;
        test_addr[2124] = 334;
        test_data[2124] = 33'd367405373;
        test_addr[2125] = 335;
        test_data[2125] = 33'd2170132500;
        test_addr[2126] = 336;
        test_data[2126] = 33'd5302575814;
        test_addr[2127] = 337;
        test_data[2127] = 33'd3038999267;
        test_addr[2128] = 338;
        test_data[2128] = 33'd4373850171;
        test_addr[2129] = 339;
        test_data[2129] = 33'd214478531;
        test_addr[2130] = 340;
        test_data[2130] = 33'd5600733017;
        test_addr[2131] = 341;
        test_data[2131] = 33'd742447467;
        test_addr[2132] = 342;
        test_data[2132] = 33'd1626249509;
        test_addr[2133] = 343;
        test_data[2133] = 33'd1398640096;
        test_addr[2134] = 991;
        test_data[2134] = 33'd961558183;
        test_addr[2135] = 992;
        test_data[2135] = 33'd7620102813;
        test_addr[2136] = 993;
        test_data[2136] = 33'd1150199168;
        test_addr[2137] = 994;
        test_data[2137] = 33'd493598879;
        test_addr[2138] = 995;
        test_data[2138] = 33'd7401391790;
        test_addr[2139] = 973;
        test_data[2139] = 33'd6493528335;
        test_addr[2140] = 974;
        test_data[2140] = 33'd2963070664;
        test_addr[2141] = 975;
        test_data[2141] = 33'd900993035;
        test_addr[2142] = 976;
        test_data[2142] = 33'd6170795515;
        test_addr[2143] = 977;
        test_data[2143] = 33'd1367094021;
        test_addr[2144] = 978;
        test_data[2144] = 33'd612406700;
        test_addr[2145] = 979;
        test_data[2145] = 33'd1047521573;
        test_addr[2146] = 980;
        test_data[2146] = 33'd3721886817;
        test_addr[2147] = 981;
        test_data[2147] = 33'd6910575997;
        test_addr[2148] = 982;
        test_data[2148] = 33'd2064422908;
        test_addr[2149] = 983;
        test_data[2149] = 33'd1240550962;
        test_addr[2150] = 984;
        test_data[2150] = 33'd7127907497;
        test_addr[2151] = 985;
        test_data[2151] = 33'd2426054176;
        test_addr[2152] = 986;
        test_data[2152] = 33'd3998934162;
        test_addr[2153] = 987;
        test_data[2153] = 33'd2162629260;
        test_addr[2154] = 996;
        test_data[2154] = 33'd103670533;
        test_addr[2155] = 997;
        test_data[2155] = 33'd5797150567;
        test_addr[2156] = 998;
        test_data[2156] = 33'd8429990815;
        test_addr[2157] = 999;
        test_data[2157] = 33'd811944595;
        test_addr[2158] = 1000;
        test_data[2158] = 33'd1407009352;
        test_addr[2159] = 1001;
        test_data[2159] = 33'd3133226956;
        test_addr[2160] = 1002;
        test_data[2160] = 33'd1816079453;
        test_addr[2161] = 1003;
        test_data[2161] = 33'd276489340;
        test_addr[2162] = 1004;
        test_data[2162] = 33'd4090172265;
        test_addr[2163] = 1005;
        test_data[2163] = 33'd1735952530;
        test_addr[2164] = 1006;
        test_data[2164] = 33'd1873145601;
        test_addr[2165] = 525;
        test_data[2165] = 33'd2372613957;
        test_addr[2166] = 526;
        test_data[2166] = 33'd6417240089;
        test_addr[2167] = 527;
        test_data[2167] = 33'd1738182943;
        test_addr[2168] = 528;
        test_data[2168] = 33'd664804818;
        test_addr[2169] = 529;
        test_data[2169] = 33'd5056814047;
        test_addr[2170] = 1007;
        test_data[2170] = 33'd635148783;
        test_addr[2171] = 1008;
        test_data[2171] = 33'd2350202510;
        test_addr[2172] = 1009;
        test_data[2172] = 33'd7990228779;
        test_addr[2173] = 1010;
        test_data[2173] = 33'd1146572673;
        test_addr[2174] = 69;
        test_data[2174] = 33'd7628867222;
        test_addr[2175] = 70;
        test_data[2175] = 33'd5031679761;
        test_addr[2176] = 71;
        test_data[2176] = 33'd7783843361;
        test_addr[2177] = 72;
        test_data[2177] = 33'd3745474962;
        test_addr[2178] = 73;
        test_data[2178] = 33'd7572833137;
        test_addr[2179] = 74;
        test_data[2179] = 33'd1195861608;
        test_addr[2180] = 75;
        test_data[2180] = 33'd3391000377;
        test_addr[2181] = 76;
        test_data[2181] = 33'd1051232611;
        test_addr[2182] = 77;
        test_data[2182] = 33'd2422841240;
        test_addr[2183] = 78;
        test_data[2183] = 33'd3591490314;
        test_addr[2184] = 79;
        test_data[2184] = 33'd466432104;
        test_addr[2185] = 80;
        test_data[2185] = 33'd3440150321;
        test_addr[2186] = 81;
        test_data[2186] = 33'd2609650108;
        test_addr[2187] = 1011;
        test_data[2187] = 33'd8201929314;
        test_addr[2188] = 1012;
        test_data[2188] = 33'd128963949;
        test_addr[2189] = 1013;
        test_data[2189] = 33'd7698810023;
        test_addr[2190] = 1014;
        test_data[2190] = 33'd7650473881;
        test_addr[2191] = 1015;
        test_data[2191] = 33'd8870532;
        test_addr[2192] = 283;
        test_data[2192] = 33'd4134955926;
        test_addr[2193] = 284;
        test_data[2193] = 33'd1470833253;
        test_addr[2194] = 285;
        test_data[2194] = 33'd5510154728;
        test_addr[2195] = 286;
        test_data[2195] = 33'd1109364526;
        test_addr[2196] = 287;
        test_data[2196] = 33'd2077233220;
        test_addr[2197] = 288;
        test_data[2197] = 33'd4027136949;
        test_addr[2198] = 289;
        test_data[2198] = 33'd940573815;
        test_addr[2199] = 290;
        test_data[2199] = 33'd7635288433;
        test_addr[2200] = 291;
        test_data[2200] = 33'd2648754452;
        test_addr[2201] = 292;
        test_data[2201] = 33'd3646512956;
        test_addr[2202] = 293;
        test_data[2202] = 33'd120765790;
        test_addr[2203] = 294;
        test_data[2203] = 33'd2357551952;
        test_addr[2204] = 1016;
        test_data[2204] = 33'd7095153347;
        test_addr[2205] = 1017;
        test_data[2205] = 33'd3197795730;
        test_addr[2206] = 1018;
        test_data[2206] = 33'd2750972131;
        test_addr[2207] = 1019;
        test_data[2207] = 33'd2061468658;
        test_addr[2208] = 1020;
        test_data[2208] = 33'd2219406155;
        test_addr[2209] = 1021;
        test_data[2209] = 33'd5546293307;
        test_addr[2210] = 1022;
        test_data[2210] = 33'd2746665182;
        test_addr[2211] = 1023;
        test_data[2211] = 33'd4086440552;
        test_addr[2212] = 0;
        test_data[2212] = 33'd5272133053;
        test_addr[2213] = 1;
        test_data[2213] = 33'd1864485560;
        test_addr[2214] = 2;
        test_data[2214] = 33'd1953611785;
        test_addr[2215] = 3;
        test_data[2215] = 33'd3350406635;
        test_addr[2216] = 4;
        test_data[2216] = 33'd1463761539;
        test_addr[2217] = 5;
        test_data[2217] = 33'd2154190107;
        test_addr[2218] = 6;
        test_data[2218] = 33'd1594182125;
        test_addr[2219] = 7;
        test_data[2219] = 33'd338412474;
        test_addr[2220] = 8;
        test_data[2220] = 33'd1742786174;
        test_addr[2221] = 9;
        test_data[2221] = 33'd6255462504;
        test_addr[2222] = 10;
        test_data[2222] = 33'd4271687727;
        test_addr[2223] = 11;
        test_data[2223] = 33'd3967754806;
        test_addr[2224] = 12;
        test_data[2224] = 33'd1768449257;
        test_addr[2225] = 13;
        test_data[2225] = 33'd4582673823;
        test_addr[2226] = 14;
        test_data[2226] = 33'd2631202414;
        test_addr[2227] = 15;
        test_data[2227] = 33'd1119003857;
        test_addr[2228] = 16;
        test_data[2228] = 33'd3925987810;
        test_addr[2229] = 17;
        test_data[2229] = 33'd7601994171;
        test_addr[2230] = 18;
        test_data[2230] = 33'd1569000094;
        test_addr[2231] = 19;
        test_data[2231] = 33'd3323511223;
        test_addr[2232] = 20;
        test_data[2232] = 33'd7763637297;
        test_addr[2233] = 21;
        test_data[2233] = 33'd1201537761;
        test_addr[2234] = 22;
        test_data[2234] = 33'd4914980157;
        test_addr[2235] = 23;
        test_data[2235] = 33'd241469200;
        test_addr[2236] = 24;
        test_data[2236] = 33'd8069725484;
        test_addr[2237] = 25;
        test_data[2237] = 33'd3473148738;
        test_addr[2238] = 236;
        test_data[2238] = 33'd5032169204;
        test_addr[2239] = 237;
        test_data[2239] = 33'd1695743965;
        test_addr[2240] = 238;
        test_data[2240] = 33'd2030143949;
        test_addr[2241] = 239;
        test_data[2241] = 33'd980297125;
        test_addr[2242] = 240;
        test_data[2242] = 33'd2785262700;
        test_addr[2243] = 26;
        test_data[2243] = 33'd3022536064;
        test_addr[2244] = 27;
        test_data[2244] = 33'd1798709310;
        test_addr[2245] = 28;
        test_data[2245] = 33'd4030679079;
        test_addr[2246] = 29;
        test_data[2246] = 33'd3629881189;
        test_addr[2247] = 30;
        test_data[2247] = 33'd7348792991;
        test_addr[2248] = 31;
        test_data[2248] = 33'd3527005491;
        test_addr[2249] = 32;
        test_data[2249] = 33'd3844512050;
        test_addr[2250] = 33;
        test_data[2250] = 33'd6220033436;
        test_addr[2251] = 34;
        test_data[2251] = 33'd4655747509;
        test_addr[2252] = 35;
        test_data[2252] = 33'd5193387947;
        test_addr[2253] = 920;
        test_data[2253] = 33'd5770974348;
        test_addr[2254] = 921;
        test_data[2254] = 33'd2992114596;
        test_addr[2255] = 922;
        test_data[2255] = 33'd6605063592;
        test_addr[2256] = 923;
        test_data[2256] = 33'd3334114139;
        test_addr[2257] = 924;
        test_data[2257] = 33'd2084629605;
        test_addr[2258] = 925;
        test_data[2258] = 33'd2610089944;
        test_addr[2259] = 926;
        test_data[2259] = 33'd3145315055;
        test_addr[2260] = 927;
        test_data[2260] = 33'd425505923;
        test_addr[2261] = 36;
        test_data[2261] = 33'd1441993322;
        test_addr[2262] = 37;
        test_data[2262] = 33'd3077452828;
        test_addr[2263] = 38;
        test_data[2263] = 33'd179744430;
        test_addr[2264] = 39;
        test_data[2264] = 33'd7004155242;
        test_addr[2265] = 40;
        test_data[2265] = 33'd710895914;
        test_addr[2266] = 41;
        test_data[2266] = 33'd2505013171;
        test_addr[2267] = 42;
        test_data[2267] = 33'd4114111253;
        test_addr[2268] = 43;
        test_data[2268] = 33'd1598694208;
        test_addr[2269] = 44;
        test_data[2269] = 33'd498645939;
        test_addr[2270] = 1014;
        test_data[2270] = 33'd3355506585;
        test_addr[2271] = 1015;
        test_data[2271] = 33'd8870532;
        test_addr[2272] = 1016;
        test_data[2272] = 33'd6089922898;
        test_addr[2273] = 1017;
        test_data[2273] = 33'd6570108758;
        test_addr[2274] = 1018;
        test_data[2274] = 33'd2750972131;
        test_addr[2275] = 1019;
        test_data[2275] = 33'd2061468658;
        test_addr[2276] = 1020;
        test_data[2276] = 33'd6106928616;
        test_addr[2277] = 1021;
        test_data[2277] = 33'd1251326011;
        test_addr[2278] = 1022;
        test_data[2278] = 33'd2746665182;
        test_addr[2279] = 1023;
        test_data[2279] = 33'd7631555268;
        test_addr[2280] = 0;
        test_data[2280] = 33'd977165757;
        test_addr[2281] = 1;
        test_data[2281] = 33'd5172932759;
        test_addr[2282] = 2;
        test_data[2282] = 33'd1953611785;
        test_addr[2283] = 3;
        test_data[2283] = 33'd3350406635;
        test_addr[2284] = 4;
        test_data[2284] = 33'd6969189185;
        test_addr[2285] = 5;
        test_data[2285] = 33'd2154190107;
        test_addr[2286] = 6;
        test_data[2286] = 33'd6081423377;
        test_addr[2287] = 7;
        test_data[2287] = 33'd338412474;
        test_addr[2288] = 8;
        test_data[2288] = 33'd1742786174;
        test_addr[2289] = 45;
        test_data[2289] = 33'd2757741745;
        test_addr[2290] = 46;
        test_data[2290] = 33'd317333202;
        test_addr[2291] = 47;
        test_data[2291] = 33'd5522597370;
        test_addr[2292] = 48;
        test_data[2292] = 33'd2577690104;
        test_addr[2293] = 49;
        test_data[2293] = 33'd7898266710;
        test_addr[2294] = 50;
        test_data[2294] = 33'd7846664864;
        test_addr[2295] = 51;
        test_data[2295] = 33'd3352351002;
        test_addr[2296] = 52;
        test_data[2296] = 33'd6484524762;
        test_addr[2297] = 53;
        test_data[2297] = 33'd2097143458;
        test_addr[2298] = 54;
        test_data[2298] = 33'd2988819932;
        test_addr[2299] = 55;
        test_data[2299] = 33'd2230608892;
        test_addr[2300] = 56;
        test_data[2300] = 33'd4190953127;
        test_addr[2301] = 57;
        test_data[2301] = 33'd2320754702;
        test_addr[2302] = 58;
        test_data[2302] = 33'd3203147784;
        test_addr[2303] = 59;
        test_data[2303] = 33'd3417772745;
        test_addr[2304] = 60;
        test_data[2304] = 33'd1830269684;
        test_addr[2305] = 10;
        test_data[2305] = 33'd4271687727;
        test_addr[2306] = 11;
        test_data[2306] = 33'd3967754806;
        test_addr[2307] = 12;
        test_data[2307] = 33'd1768449257;
        test_addr[2308] = 13;
        test_data[2308] = 33'd4830922811;
        test_addr[2309] = 14;
        test_data[2309] = 33'd5126967643;
        test_addr[2310] = 61;
        test_data[2310] = 33'd2209095858;
        test_addr[2311] = 324;
        test_data[2311] = 33'd2439471225;
        test_addr[2312] = 325;
        test_data[2312] = 33'd8099382805;
        test_addr[2313] = 326;
        test_data[2313] = 33'd8185249838;
        test_addr[2314] = 327;
        test_data[2314] = 33'd318989378;
        test_addr[2315] = 328;
        test_data[2315] = 33'd3131202390;
        test_addr[2316] = 329;
        test_data[2316] = 33'd3139848229;
        test_addr[2317] = 330;
        test_data[2317] = 33'd5126305773;
        test_addr[2318] = 331;
        test_data[2318] = 33'd2887064224;
        test_addr[2319] = 332;
        test_data[2319] = 33'd2382769822;
        test_addr[2320] = 333;
        test_data[2320] = 33'd1462324255;
        test_addr[2321] = 62;
        test_data[2321] = 33'd504570280;
        test_addr[2322] = 63;
        test_data[2322] = 33'd4143158891;
        test_addr[2323] = 64;
        test_data[2323] = 33'd1705434463;
        test_addr[2324] = 65;
        test_data[2324] = 33'd6955468322;
        test_addr[2325] = 66;
        test_data[2325] = 33'd7969941461;
        test_addr[2326] = 67;
        test_data[2326] = 33'd2781999553;
        test_addr[2327] = 68;
        test_data[2327] = 33'd7211945344;
        test_addr[2328] = 69;
        test_data[2328] = 33'd3333899926;
        test_addr[2329] = 70;
        test_data[2329] = 33'd736712465;
        test_addr[2330] = 71;
        test_data[2330] = 33'd6151953823;
        test_addr[2331] = 33;
        test_data[2331] = 33'd1925066140;
        test_addr[2332] = 34;
        test_data[2332] = 33'd360780213;
        test_addr[2333] = 35;
        test_data[2333] = 33'd898420651;
        test_addr[2334] = 36;
        test_data[2334] = 33'd7523352331;
        test_addr[2335] = 37;
        test_data[2335] = 33'd3077452828;
        test_addr[2336] = 72;
        test_data[2336] = 33'd3745474962;
        test_addr[2337] = 73;
        test_data[2337] = 33'd3277865841;
        test_addr[2338] = 74;
        test_data[2338] = 33'd1195861608;
        test_addr[2339] = 75;
        test_data[2339] = 33'd3391000377;
        test_addr[2340] = 76;
        test_data[2340] = 33'd1051232611;
        test_addr[2341] = 77;
        test_data[2341] = 33'd2422841240;
        test_addr[2342] = 78;
        test_data[2342] = 33'd3591490314;
        test_addr[2343] = 79;
        test_data[2343] = 33'd4648328243;
        test_addr[2344] = 80;
        test_data[2344] = 33'd3440150321;
        test_addr[2345] = 81;
        test_data[2345] = 33'd2609650108;
        test_addr[2346] = 82;
        test_data[2346] = 33'd1149693843;
        test_addr[2347] = 83;
        test_data[2347] = 33'd176121797;
        test_addr[2348] = 728;
        test_data[2348] = 33'd1284317235;
        test_addr[2349] = 729;
        test_data[2349] = 33'd919345546;
        test_addr[2350] = 730;
        test_data[2350] = 33'd4067928788;
        test_addr[2351] = 731;
        test_data[2351] = 33'd1353510671;
        test_addr[2352] = 732;
        test_data[2352] = 33'd6000833766;
        test_addr[2353] = 733;
        test_data[2353] = 33'd8165455448;
        test_addr[2354] = 734;
        test_data[2354] = 33'd4496695338;
        test_addr[2355] = 735;
        test_data[2355] = 33'd6265892489;
        test_addr[2356] = 736;
        test_data[2356] = 33'd2719855705;
        test_addr[2357] = 737;
        test_data[2357] = 33'd7442161535;
        test_addr[2358] = 84;
        test_data[2358] = 33'd5443080443;
        test_addr[2359] = 85;
        test_data[2359] = 33'd3382751907;
        test_addr[2360] = 86;
        test_data[2360] = 33'd623629618;
        test_addr[2361] = 87;
        test_data[2361] = 33'd3303907992;
        test_addr[2362] = 88;
        test_data[2362] = 33'd5906344003;
        test_addr[2363] = 89;
        test_data[2363] = 33'd1036241526;
        test_addr[2364] = 90;
        test_data[2364] = 33'd548807498;
        test_addr[2365] = 91;
        test_data[2365] = 33'd4425844943;
        test_addr[2366] = 92;
        test_data[2366] = 33'd6570401415;
        test_addr[2367] = 204;
        test_data[2367] = 33'd3073370316;
        test_addr[2368] = 205;
        test_data[2368] = 33'd6832772999;
        test_addr[2369] = 206;
        test_data[2369] = 33'd871555750;
        test_addr[2370] = 93;
        test_data[2370] = 33'd284207449;
        test_addr[2371] = 94;
        test_data[2371] = 33'd4015470161;
        test_addr[2372] = 95;
        test_data[2372] = 33'd6645332227;
        test_addr[2373] = 96;
        test_data[2373] = 33'd1425630043;
        test_addr[2374] = 97;
        test_data[2374] = 33'd3179244300;
        test_addr[2375] = 98;
        test_data[2375] = 33'd4401623969;
        test_addr[2376] = 99;
        test_data[2376] = 33'd6083966729;
        test_addr[2377] = 877;
        test_data[2377] = 33'd2926156055;
        test_addr[2378] = 878;
        test_data[2378] = 33'd3725508185;
        test_addr[2379] = 879;
        test_data[2379] = 33'd6284484629;
        test_addr[2380] = 880;
        test_data[2380] = 33'd3264573792;
        test_addr[2381] = 881;
        test_data[2381] = 33'd156207808;
        test_addr[2382] = 882;
        test_data[2382] = 33'd3569824834;
        test_addr[2383] = 883;
        test_data[2383] = 33'd6200842172;
        test_addr[2384] = 884;
        test_data[2384] = 33'd7485881606;
        test_addr[2385] = 885;
        test_data[2385] = 33'd3458389258;
        test_addr[2386] = 886;
        test_data[2386] = 33'd4811166535;
        test_addr[2387] = 887;
        test_data[2387] = 33'd2507313658;
        test_addr[2388] = 888;
        test_data[2388] = 33'd397640837;
        test_addr[2389] = 889;
        test_data[2389] = 33'd1528309135;
        test_addr[2390] = 890;
        test_data[2390] = 33'd7699099764;
        test_addr[2391] = 891;
        test_data[2391] = 33'd7756056860;
        test_addr[2392] = 892;
        test_data[2392] = 33'd8421272827;
        test_addr[2393] = 893;
        test_data[2393] = 33'd177830993;
        test_addr[2394] = 100;
        test_data[2394] = 33'd1558129631;
        test_addr[2395] = 101;
        test_data[2395] = 33'd2188618610;
        test_addr[2396] = 102;
        test_data[2396] = 33'd3632082374;
        test_addr[2397] = 103;
        test_data[2397] = 33'd2907570000;
        test_addr[2398] = 104;
        test_data[2398] = 33'd2404063296;
        test_addr[2399] = 105;
        test_data[2399] = 33'd1914703890;
        test_addr[2400] = 106;
        test_data[2400] = 33'd568746040;
        test_addr[2401] = 107;
        test_data[2401] = 33'd2329785644;
        test_addr[2402] = 652;
        test_data[2402] = 33'd3998291136;
        test_addr[2403] = 653;
        test_data[2403] = 33'd8036140886;
        test_addr[2404] = 108;
        test_data[2404] = 33'd8154949647;
        test_addr[2405] = 109;
        test_data[2405] = 33'd2828290416;
        test_addr[2406] = 110;
        test_data[2406] = 33'd3917257109;
        test_addr[2407] = 111;
        test_data[2407] = 33'd4583562168;
        test_addr[2408] = 112;
        test_data[2408] = 33'd1611235687;
        test_addr[2409] = 113;
        test_data[2409] = 33'd3918457011;
        test_addr[2410] = 114;
        test_data[2410] = 33'd5028372430;
        test_addr[2411] = 115;
        test_data[2411] = 33'd4585425408;
        test_addr[2412] = 159;
        test_data[2412] = 33'd8009700248;
        test_addr[2413] = 160;
        test_data[2413] = 33'd2220794859;
        test_addr[2414] = 116;
        test_data[2414] = 33'd1148833960;
        test_addr[2415] = 117;
        test_data[2415] = 33'd2672303755;
        test_addr[2416] = 903;
        test_data[2416] = 33'd486481265;
        test_addr[2417] = 904;
        test_data[2417] = 33'd299855562;
        test_addr[2418] = 905;
        test_data[2418] = 33'd8089781019;
        test_addr[2419] = 906;
        test_data[2419] = 33'd7430002691;
        test_addr[2420] = 907;
        test_data[2420] = 33'd1829404985;
        test_addr[2421] = 908;
        test_data[2421] = 33'd6130930004;
        test_addr[2422] = 909;
        test_data[2422] = 33'd4647221617;
        test_addr[2423] = 910;
        test_data[2423] = 33'd5927051762;
        test_addr[2424] = 911;
        test_data[2424] = 33'd806648968;
        test_addr[2425] = 912;
        test_data[2425] = 33'd4686496519;
        test_addr[2426] = 118;
        test_data[2426] = 33'd7352648691;
        test_addr[2427] = 340;
        test_data[2427] = 33'd7631007457;
        test_addr[2428] = 341;
        test_data[2428] = 33'd742447467;
        test_addr[2429] = 342;
        test_data[2429] = 33'd1626249509;
        test_addr[2430] = 343;
        test_data[2430] = 33'd1398640096;
        test_addr[2431] = 344;
        test_data[2431] = 33'd281373290;
        test_addr[2432] = 345;
        test_data[2432] = 33'd7335172044;
        test_addr[2433] = 346;
        test_data[2433] = 33'd571024672;
        test_addr[2434] = 347;
        test_data[2434] = 33'd6940813752;
        test_addr[2435] = 348;
        test_data[2435] = 33'd3632034653;
        test_addr[2436] = 349;
        test_data[2436] = 33'd516820221;
        test_addr[2437] = 119;
        test_data[2437] = 33'd8586247483;
        test_addr[2438] = 120;
        test_data[2438] = 33'd4983909213;
        test_addr[2439] = 121;
        test_data[2439] = 33'd5279619265;
        test_addr[2440] = 122;
        test_data[2440] = 33'd1367201542;
        test_addr[2441] = 123;
        test_data[2441] = 33'd313859363;
        test_addr[2442] = 124;
        test_data[2442] = 33'd8041912983;
        test_addr[2443] = 125;
        test_data[2443] = 33'd1825838587;
        test_addr[2444] = 126;
        test_data[2444] = 33'd4377020472;
        test_addr[2445] = 127;
        test_data[2445] = 33'd6863717041;
        test_addr[2446] = 128;
        test_data[2446] = 33'd2661708367;
        test_addr[2447] = 129;
        test_data[2447] = 33'd4838522692;
        test_addr[2448] = 130;
        test_data[2448] = 33'd454112648;
        test_addr[2449] = 98;
        test_data[2449] = 33'd106656673;
        test_addr[2450] = 99;
        test_data[2450] = 33'd1788999433;
        test_addr[2451] = 100;
        test_data[2451] = 33'd7661181908;
        test_addr[2452] = 131;
        test_data[2452] = 33'd5199504147;
        test_addr[2453] = 132;
        test_data[2453] = 33'd7675725971;
        test_addr[2454] = 133;
        test_data[2454] = 33'd1549772363;
        test_addr[2455] = 134;
        test_data[2455] = 33'd2986512865;
        test_addr[2456] = 135;
        test_data[2456] = 33'd1960021159;
        test_addr[2457] = 136;
        test_data[2457] = 33'd8552008386;
        test_addr[2458] = 137;
        test_data[2458] = 33'd4030908906;
        test_addr[2459] = 138;
        test_data[2459] = 33'd2117276309;
        test_addr[2460] = 139;
        test_data[2460] = 33'd643785746;
        test_addr[2461] = 140;
        test_data[2461] = 33'd6630848110;
        test_addr[2462] = 141;
        test_data[2462] = 33'd3385276041;
        test_addr[2463] = 142;
        test_data[2463] = 33'd2889759130;
        test_addr[2464] = 143;
        test_data[2464] = 33'd7456523381;
        test_addr[2465] = 144;
        test_data[2465] = 33'd3584443635;
        test_addr[2466] = 145;
        test_data[2466] = 33'd2276121759;
        test_addr[2467] = 146;
        test_data[2467] = 33'd1978812597;
        test_addr[2468] = 147;
        test_data[2468] = 33'd3498313420;
        test_addr[2469] = 148;
        test_data[2469] = 33'd4014633640;
        test_addr[2470] = 149;
        test_data[2470] = 33'd5347881512;
        test_addr[2471] = 6;
        test_data[2471] = 33'd1786456081;
        test_addr[2472] = 7;
        test_data[2472] = 33'd6230351071;
        test_addr[2473] = 8;
        test_data[2473] = 33'd7723818367;
        test_addr[2474] = 9;
        test_data[2474] = 33'd1960495208;
        test_addr[2475] = 10;
        test_data[2475] = 33'd4271687727;
        test_addr[2476] = 11;
        test_data[2476] = 33'd7939535672;
        test_addr[2477] = 12;
        test_data[2477] = 33'd1768449257;
        test_addr[2478] = 13;
        test_data[2478] = 33'd535955515;
        test_addr[2479] = 14;
        test_data[2479] = 33'd832000347;
        test_addr[2480] = 15;
        test_data[2480] = 33'd1119003857;
        test_addr[2481] = 16;
        test_data[2481] = 33'd3925987810;
        test_addr[2482] = 17;
        test_data[2482] = 33'd3307026875;
        test_addr[2483] = 18;
        test_data[2483] = 33'd1569000094;
        test_addr[2484] = 150;
        test_data[2484] = 33'd1729930243;
        test_addr[2485] = 151;
        test_data[2485] = 33'd6885124379;
        test_addr[2486] = 152;
        test_data[2486] = 33'd6602432073;
        test_addr[2487] = 153;
        test_data[2487] = 33'd352254805;
        test_addr[2488] = 154;
        test_data[2488] = 33'd8377983174;
        test_addr[2489] = 155;
        test_data[2489] = 33'd6217604989;
        test_addr[2490] = 156;
        test_data[2490] = 33'd1324821377;
        test_addr[2491] = 157;
        test_data[2491] = 33'd2090366039;
        test_addr[2492] = 158;
        test_data[2492] = 33'd5456442795;
        test_addr[2493] = 159;
        test_data[2493] = 33'd5898995500;
        test_addr[2494] = 160;
        test_data[2494] = 33'd2220794859;
        test_addr[2495] = 161;
        test_data[2495] = 33'd3906768938;
        test_addr[2496] = 162;
        test_data[2496] = 33'd775522268;
        test_addr[2497] = 163;
        test_data[2497] = 33'd8509088075;
        test_addr[2498] = 164;
        test_data[2498] = 33'd2460820341;
        test_addr[2499] = 165;
        test_data[2499] = 33'd6082145369;
        test_addr[2500] = 166;
        test_data[2500] = 33'd7002908252;
        test_addr[2501] = 167;
        test_data[2501] = 33'd1936248238;
        test_addr[2502] = 168;
        test_data[2502] = 33'd6273700389;
        test_addr[2503] = 169;
        test_data[2503] = 33'd2652621613;
        test_addr[2504] = 170;
        test_data[2504] = 33'd5199623728;
        test_addr[2505] = 171;
        test_data[2505] = 33'd3511614128;
        test_addr[2506] = 172;
        test_data[2506] = 33'd4198004977;
        test_addr[2507] = 173;
        test_data[2507] = 33'd4797826549;
        test_addr[2508] = 988;
        test_data[2508] = 33'd1189533474;
        test_addr[2509] = 989;
        test_data[2509] = 33'd6915543312;
        test_addr[2510] = 174;
        test_data[2510] = 33'd2285112422;
        test_addr[2511] = 175;
        test_data[2511] = 33'd3567745488;
        test_addr[2512] = 176;
        test_data[2512] = 33'd2422858599;
        test_addr[2513] = 177;
        test_data[2513] = 33'd4649219896;
        test_addr[2514] = 178;
        test_data[2514] = 33'd745299376;
        test_addr[2515] = 179;
        test_data[2515] = 33'd6714553003;
        test_addr[2516] = 180;
        test_data[2516] = 33'd4240384840;
        test_addr[2517] = 181;
        test_data[2517] = 33'd2156248305;
        test_addr[2518] = 182;
        test_data[2518] = 33'd1222529405;
        test_addr[2519] = 183;
        test_data[2519] = 33'd4192569996;
        test_addr[2520] = 184;
        test_data[2520] = 33'd8535355262;
        test_addr[2521] = 185;
        test_data[2521] = 33'd8159830687;
        test_addr[2522] = 186;
        test_data[2522] = 33'd2175561490;
        test_addr[2523] = 187;
        test_data[2523] = 33'd4277874876;
        test_addr[2524] = 188;
        test_data[2524] = 33'd128496091;
        test_addr[2525] = 189;
        test_data[2525] = 33'd133639369;
        test_addr[2526] = 190;
        test_data[2526] = 33'd6313215124;
        test_addr[2527] = 191;
        test_data[2527] = 33'd8246956740;
        test_addr[2528] = 192;
        test_data[2528] = 33'd275041321;
        test_addr[2529] = 193;
        test_data[2529] = 33'd5943030237;
        test_addr[2530] = 194;
        test_data[2530] = 33'd6512977942;
        test_addr[2531] = 971;
        test_data[2531] = 33'd5945151923;
        test_addr[2532] = 972;
        test_data[2532] = 33'd2381619306;
        test_addr[2533] = 973;
        test_data[2533] = 33'd2198561039;
        test_addr[2534] = 974;
        test_data[2534] = 33'd8200593194;
        test_addr[2535] = 195;
        test_data[2535] = 33'd3241511229;
        test_addr[2536] = 196;
        test_data[2536] = 33'd1811402878;
        test_addr[2537] = 197;
        test_data[2537] = 33'd7221533045;
        test_addr[2538] = 804;
        test_data[2538] = 33'd7052923694;
        test_addr[2539] = 805;
        test_data[2539] = 33'd5880258990;
        test_addr[2540] = 806;
        test_data[2540] = 33'd1359101487;
        test_addr[2541] = 807;
        test_data[2541] = 33'd540490609;
        test_addr[2542] = 808;
        test_data[2542] = 33'd4179863201;
        test_addr[2543] = 809;
        test_data[2543] = 33'd3766935983;
        test_addr[2544] = 810;
        test_data[2544] = 33'd4828242253;
        test_addr[2545] = 811;
        test_data[2545] = 33'd5013471150;
        test_addr[2546] = 812;
        test_data[2546] = 33'd6342945479;
        test_addr[2547] = 198;
        test_data[2547] = 33'd1771443269;
        test_addr[2548] = 199;
        test_data[2548] = 33'd285609981;
        test_addr[2549] = 200;
        test_data[2549] = 33'd5909894956;
        test_addr[2550] = 201;
        test_data[2550] = 33'd4682522543;
        test_addr[2551] = 980;
        test_data[2551] = 33'd5196539160;
        test_addr[2552] = 981;
        test_data[2552] = 33'd7010175952;
        test_addr[2553] = 982;
        test_data[2553] = 33'd2064422908;
        test_addr[2554] = 983;
        test_data[2554] = 33'd1240550962;
        test_addr[2555] = 984;
        test_data[2555] = 33'd5811921495;
        test_addr[2556] = 985;
        test_data[2556] = 33'd2426054176;
        test_addr[2557] = 986;
        test_data[2557] = 33'd3998934162;
        test_addr[2558] = 987;
        test_data[2558] = 33'd2162629260;
        test_addr[2559] = 988;
        test_data[2559] = 33'd6708303644;
        test_addr[2560] = 989;
        test_data[2560] = 33'd2620576016;
        test_addr[2561] = 990;
        test_data[2561] = 33'd431413773;
        test_addr[2562] = 202;
        test_data[2562] = 33'd6921128689;
        test_addr[2563] = 203;
        test_data[2563] = 33'd1663091370;
        test_addr[2564] = 204;
        test_data[2564] = 33'd7752091514;
        test_addr[2565] = 205;
        test_data[2565] = 33'd2537805703;
        test_addr[2566] = 206;
        test_data[2566] = 33'd871555750;
        test_addr[2567] = 207;
        test_data[2567] = 33'd3823761644;
        test_addr[2568] = 208;
        test_data[2568] = 33'd3010632164;
        test_addr[2569] = 288;
        test_data[2569] = 33'd7066161205;
        test_addr[2570] = 289;
        test_data[2570] = 33'd940573815;
        test_addr[2571] = 290;
        test_data[2571] = 33'd6774055835;
        test_addr[2572] = 291;
        test_data[2572] = 33'd2648754452;
        test_addr[2573] = 209;
        test_data[2573] = 33'd7202450869;
        test_addr[2574] = 210;
        test_data[2574] = 33'd391446383;
        test_addr[2575] = 900;
        test_data[2575] = 33'd2081706384;
        test_addr[2576] = 901;
        test_data[2576] = 33'd1604865859;
        test_addr[2577] = 902;
        test_data[2577] = 33'd3762112714;
        test_addr[2578] = 903;
        test_data[2578] = 33'd486481265;
        test_addr[2579] = 904;
        test_data[2579] = 33'd299855562;
        test_addr[2580] = 905;
        test_data[2580] = 33'd3794813723;
        test_addr[2581] = 906;
        test_data[2581] = 33'd3135035395;
        test_addr[2582] = 907;
        test_data[2582] = 33'd1829404985;
        test_addr[2583] = 908;
        test_data[2583] = 33'd1835962708;
        test_addr[2584] = 211;
        test_data[2584] = 33'd7044103130;
        test_addr[2585] = 212;
        test_data[2585] = 33'd7742942298;
        test_addr[2586] = 213;
        test_data[2586] = 33'd8489706716;
        test_addr[2587] = 214;
        test_data[2587] = 33'd4759522780;
        test_addr[2588] = 215;
        test_data[2588] = 33'd4957648746;
        test_addr[2589] = 216;
        test_data[2589] = 33'd708341535;
        test_addr[2590] = 217;
        test_data[2590] = 33'd7597289486;
        test_addr[2591] = 218;
        test_data[2591] = 33'd1182784850;
        test_addr[2592] = 219;
        test_data[2592] = 33'd2689063963;
        test_addr[2593] = 888;
        test_data[2593] = 33'd7377037149;
        test_addr[2594] = 889;
        test_data[2594] = 33'd5910934898;
        test_addr[2595] = 890;
        test_data[2595] = 33'd3404132468;
        test_addr[2596] = 891;
        test_data[2596] = 33'd3461089564;
        test_addr[2597] = 892;
        test_data[2597] = 33'd6532726900;
        test_addr[2598] = 893;
        test_data[2598] = 33'd177830993;
        test_addr[2599] = 220;
        test_data[2599] = 33'd8373386745;
        test_addr[2600] = 221;
        test_data[2600] = 33'd7528151048;
        test_addr[2601] = 222;
        test_data[2601] = 33'd4794926573;
        test_addr[2602] = 223;
        test_data[2602] = 33'd7225472110;
        test_addr[2603] = 224;
        test_data[2603] = 33'd3332430587;
        test_addr[2604] = 225;
        test_data[2604] = 33'd206097148;
        test_addr[2605] = 226;
        test_data[2605] = 33'd2883781805;
        test_addr[2606] = 227;
        test_data[2606] = 33'd5000662689;
        test_addr[2607] = 228;
        test_data[2607] = 33'd5034371648;
        test_addr[2608] = 229;
        test_data[2608] = 33'd845232644;
        test_addr[2609] = 230;
        test_data[2609] = 33'd435407810;
        test_addr[2610] = 231;
        test_data[2610] = 33'd164270080;
        test_addr[2611] = 232;
        test_data[2611] = 33'd6457463073;
        test_addr[2612] = 233;
        test_data[2612] = 33'd2304627638;
        test_addr[2613] = 234;
        test_data[2613] = 33'd2711743575;
        test_addr[2614] = 235;
        test_data[2614] = 33'd1995153683;
        test_addr[2615] = 236;
        test_data[2615] = 33'd737201908;
        test_addr[2616] = 237;
        test_data[2616] = 33'd1695743965;
        test_addr[2617] = 238;
        test_data[2617] = 33'd2030143949;
        test_addr[2618] = 239;
        test_data[2618] = 33'd980297125;
        test_addr[2619] = 240;
        test_data[2619] = 33'd5859139615;
        test_addr[2620] = 241;
        test_data[2620] = 33'd3647911902;
        test_addr[2621] = 218;
        test_data[2621] = 33'd7340064211;
        test_addr[2622] = 219;
        test_data[2622] = 33'd2689063963;
        test_addr[2623] = 220;
        test_data[2623] = 33'd7852856989;
        test_addr[2624] = 221;
        test_data[2624] = 33'd4534161241;
        test_addr[2625] = 222;
        test_data[2625] = 33'd499959277;
        test_addr[2626] = 242;
        test_data[2626] = 33'd1066521417;
        test_addr[2627] = 243;
        test_data[2627] = 33'd6892698721;
        test_addr[2628] = 244;
        test_data[2628] = 33'd2896346636;
        test_addr[2629] = 245;
        test_data[2629] = 33'd2801824671;
        test_addr[2630] = 246;
        test_data[2630] = 33'd7837856130;
        test_addr[2631] = 247;
        test_data[2631] = 33'd2088915050;
        test_addr[2632] = 248;
        test_data[2632] = 33'd7741058444;
        test_addr[2633] = 249;
        test_data[2633] = 33'd634363534;
        test_addr[2634] = 250;
        test_data[2634] = 33'd3563604010;
        test_addr[2635] = 952;
        test_data[2635] = 33'd1791314849;
        test_addr[2636] = 953;
        test_data[2636] = 33'd2693867941;
        test_addr[2637] = 954;
        test_data[2637] = 33'd2796648127;
        test_addr[2638] = 955;
        test_data[2638] = 33'd905894982;
        test_addr[2639] = 956;
        test_data[2639] = 33'd90020364;
        test_addr[2640] = 957;
        test_data[2640] = 33'd2991872276;
        test_addr[2641] = 958;
        test_data[2641] = 33'd3447221745;
        test_addr[2642] = 959;
        test_data[2642] = 33'd3794599805;
        test_addr[2643] = 960;
        test_data[2643] = 33'd3344962385;
        test_addr[2644] = 961;
        test_data[2644] = 33'd4559298786;
        test_addr[2645] = 962;
        test_data[2645] = 33'd2567179456;
        test_addr[2646] = 963;
        test_data[2646] = 33'd8457779625;
        test_addr[2647] = 251;
        test_data[2647] = 33'd7008018092;
        test_addr[2648] = 927;
        test_data[2648] = 33'd6417802278;
        test_addr[2649] = 252;
        test_data[2649] = 33'd3233104755;
        test_addr[2650] = 505;
        test_data[2650] = 33'd1706057765;
        test_addr[2651] = 506;
        test_data[2651] = 33'd847909313;
        test_addr[2652] = 507;
        test_data[2652] = 33'd7478178644;
        test_addr[2653] = 253;
        test_data[2653] = 33'd2251486923;
        test_addr[2654] = 254;
        test_data[2654] = 33'd4863868379;
        test_addr[2655] = 255;
        test_data[2655] = 33'd1613786967;
        test_addr[2656] = 256;
        test_data[2656] = 33'd3353620761;
        test_addr[2657] = 257;
        test_data[2657] = 33'd5783401445;
        test_addr[2658] = 258;
        test_data[2658] = 33'd3768261454;
        test_addr[2659] = 773;
        test_data[2659] = 33'd7114841289;
        test_addr[2660] = 774;
        test_data[2660] = 33'd9534195;
        test_addr[2661] = 775;
        test_data[2661] = 33'd7323266348;
        test_addr[2662] = 259;
        test_data[2662] = 33'd1403616719;
        test_addr[2663] = 383;
        test_data[2663] = 33'd6963298775;
        test_addr[2664] = 384;
        test_data[2664] = 33'd8174167570;
        test_addr[2665] = 385;
        test_data[2665] = 33'd5753802877;
        test_addr[2666] = 386;
        test_data[2666] = 33'd5916370253;
        test_addr[2667] = 387;
        test_data[2667] = 33'd6491283755;
        test_addr[2668] = 388;
        test_data[2668] = 33'd2217298716;
        test_addr[2669] = 389;
        test_data[2669] = 33'd4986008991;
        test_addr[2670] = 390;
        test_data[2670] = 33'd3947964093;
        test_addr[2671] = 391;
        test_data[2671] = 33'd4156755592;
        test_addr[2672] = 392;
        test_data[2672] = 33'd7964693986;
        test_addr[2673] = 393;
        test_data[2673] = 33'd3584816215;
        test_addr[2674] = 394;
        test_data[2674] = 33'd2343163130;
        test_addr[2675] = 395;
        test_data[2675] = 33'd3549743356;
        test_addr[2676] = 260;
        test_data[2676] = 33'd2209658087;
        test_addr[2677] = 261;
        test_data[2677] = 33'd2908678289;
        test_addr[2678] = 262;
        test_data[2678] = 33'd3668048787;
        test_addr[2679] = 263;
        test_data[2679] = 33'd5760665546;
        test_addr[2680] = 264;
        test_data[2680] = 33'd6623879302;
        test_addr[2681] = 265;
        test_data[2681] = 33'd5795405298;
        test_addr[2682] = 266;
        test_data[2682] = 33'd6655574761;
        test_addr[2683] = 267;
        test_data[2683] = 33'd5507743838;
        test_addr[2684] = 268;
        test_data[2684] = 33'd458908171;
        test_addr[2685] = 269;
        test_data[2685] = 33'd123635395;
        test_addr[2686] = 270;
        test_data[2686] = 33'd2703615357;
        test_addr[2687] = 195;
        test_data[2687] = 33'd3241511229;
        test_addr[2688] = 196;
        test_data[2688] = 33'd1811402878;
        test_addr[2689] = 197;
        test_data[2689] = 33'd2926565749;
        test_addr[2690] = 198;
        test_data[2690] = 33'd1771443269;
        test_addr[2691] = 199;
        test_data[2691] = 33'd4583338188;
        test_addr[2692] = 200;
        test_data[2692] = 33'd1614927660;
        test_addr[2693] = 201;
        test_data[2693] = 33'd387555247;
        test_addr[2694] = 202;
        test_data[2694] = 33'd2626161393;
        test_addr[2695] = 203;
        test_data[2695] = 33'd1663091370;
        test_addr[2696] = 204;
        test_data[2696] = 33'd3457124218;
        test_addr[2697] = 205;
        test_data[2697] = 33'd2537805703;
        test_addr[2698] = 271;
        test_data[2698] = 33'd4007140997;
        test_addr[2699] = 272;
        test_data[2699] = 33'd495494873;
        test_addr[2700] = 273;
        test_data[2700] = 33'd1263813313;
        test_addr[2701] = 274;
        test_data[2701] = 33'd1474849930;
        test_addr[2702] = 36;
        test_data[2702] = 33'd3228385035;
        test_addr[2703] = 37;
        test_data[2703] = 33'd3077452828;
        test_addr[2704] = 38;
        test_data[2704] = 33'd7406271556;
        test_addr[2705] = 39;
        test_data[2705] = 33'd2709187946;
        test_addr[2706] = 40;
        test_data[2706] = 33'd710895914;
        test_addr[2707] = 41;
        test_data[2707] = 33'd2505013171;
        test_addr[2708] = 42;
        test_data[2708] = 33'd4114111253;
        test_addr[2709] = 43;
        test_data[2709] = 33'd1598694208;
        test_addr[2710] = 44;
        test_data[2710] = 33'd7878506478;
        test_addr[2711] = 275;
        test_data[2711] = 33'd94646178;
        test_addr[2712] = 276;
        test_data[2712] = 33'd3369498205;
        test_addr[2713] = 277;
        test_data[2713] = 33'd76492403;
        test_addr[2714] = 278;
        test_data[2714] = 33'd3484772131;
        test_addr[2715] = 760;
        test_data[2715] = 33'd5468052640;
        test_addr[2716] = 761;
        test_data[2716] = 33'd8171783895;
        test_addr[2717] = 762;
        test_data[2717] = 33'd3993692466;
        test_addr[2718] = 763;
        test_data[2718] = 33'd930239523;
        test_addr[2719] = 279;
        test_data[2719] = 33'd1301179723;
        test_addr[2720] = 280;
        test_data[2720] = 33'd535207050;
        test_addr[2721] = 281;
        test_data[2721] = 33'd3105421778;
        test_addr[2722] = 282;
        test_data[2722] = 33'd1396158732;
        test_addr[2723] = 283;
        test_data[2723] = 33'd6024137186;
        test_addr[2724] = 284;
        test_data[2724] = 33'd1470833253;
        test_addr[2725] = 285;
        test_data[2725] = 33'd5142073086;
        test_addr[2726] = 286;
        test_data[2726] = 33'd1109364526;
        test_addr[2727] = 287;
        test_data[2727] = 33'd2077233220;
        test_addr[2728] = 288;
        test_data[2728] = 33'd2771193909;
        test_addr[2729] = 289;
        test_data[2729] = 33'd7652457687;
        test_addr[2730] = 290;
        test_data[2730] = 33'd5816581402;
        test_addr[2731] = 291;
        test_data[2731] = 33'd2648754452;
        test_addr[2732] = 292;
        test_data[2732] = 33'd8144763376;
        test_addr[2733] = 293;
        test_data[2733] = 33'd120765790;
        test_addr[2734] = 294;
        test_data[2734] = 33'd2357551952;
        test_addr[2735] = 295;
        test_data[2735] = 33'd431105951;
        test_addr[2736] = 296;
        test_data[2736] = 33'd6281365586;
        test_addr[2737] = 297;
        test_data[2737] = 33'd3193633458;
        test_addr[2738] = 298;
        test_data[2738] = 33'd6297611830;
        test_addr[2739] = 299;
        test_data[2739] = 33'd6458166644;
        test_addr[2740] = 300;
        test_data[2740] = 33'd1880021582;
        test_addr[2741] = 301;
        test_data[2741] = 33'd6177302279;
        test_addr[2742] = 302;
        test_data[2742] = 33'd5715156921;
        test_addr[2743] = 303;
        test_data[2743] = 33'd5573843424;
        test_addr[2744] = 304;
        test_data[2744] = 33'd460827716;
        test_addr[2745] = 305;
        test_data[2745] = 33'd1866235150;
        test_addr[2746] = 306;
        test_data[2746] = 33'd1400119106;
        test_addr[2747] = 307;
        test_data[2747] = 33'd4821889301;
        test_addr[2748] = 308;
        test_data[2748] = 33'd2611705428;
        test_addr[2749] = 309;
        test_data[2749] = 33'd3941608837;
        test_addr[2750] = 310;
        test_data[2750] = 33'd3094631771;
        test_addr[2751] = 311;
        test_data[2751] = 33'd4590676607;
        test_addr[2752] = 312;
        test_data[2752] = 33'd240548675;
        test_addr[2753] = 313;
        test_data[2753] = 33'd3069166694;
        test_addr[2754] = 314;
        test_data[2754] = 33'd2141065806;
        test_addr[2755] = 315;
        test_data[2755] = 33'd3309303920;
        test_addr[2756] = 316;
        test_data[2756] = 33'd2758457540;
        test_addr[2757] = 317;
        test_data[2757] = 33'd4112356272;
        test_addr[2758] = 338;
        test_data[2758] = 33'd78882875;
        test_addr[2759] = 339;
        test_data[2759] = 33'd214478531;
        test_addr[2760] = 340;
        test_data[2760] = 33'd3336040161;
        test_addr[2761] = 341;
        test_data[2761] = 33'd742447467;
        test_addr[2762] = 318;
        test_data[2762] = 33'd5526052598;
        test_addr[2763] = 319;
        test_data[2763] = 33'd398366425;
        test_addr[2764] = 320;
        test_data[2764] = 33'd2213105581;
        test_addr[2765] = 321;
        test_data[2765] = 33'd4078285937;
        test_addr[2766] = 322;
        test_data[2766] = 33'd5004635942;
        test_addr[2767] = 323;
        test_data[2767] = 33'd2407757486;
        test_addr[2768] = 324;
        test_data[2768] = 33'd2439471225;
        test_addr[2769] = 325;
        test_data[2769] = 33'd8229996868;
        test_addr[2770] = 326;
        test_data[2770] = 33'd7974813783;
        test_addr[2771] = 327;
        test_data[2771] = 33'd318989378;
        test_addr[2772] = 328;
        test_data[2772] = 33'd3131202390;
        test_addr[2773] = 329;
        test_data[2773] = 33'd7670674182;
        test_addr[2774] = 330;
        test_data[2774] = 33'd4456503884;
        test_addr[2775] = 331;
        test_data[2775] = 33'd2887064224;
        test_addr[2776] = 332;
        test_data[2776] = 33'd2382769822;
        test_addr[2777] = 333;
        test_data[2777] = 33'd1462324255;
        test_addr[2778] = 334;
        test_data[2778] = 33'd6177998017;
        test_addr[2779] = 335;
        test_data[2779] = 33'd2170132500;
        test_addr[2780] = 336;
        test_data[2780] = 33'd1007608518;
        test_addr[2781] = 337;
        test_data[2781] = 33'd7275875051;
        test_addr[2782] = 184;
        test_data[2782] = 33'd4240387966;
        test_addr[2783] = 185;
        test_data[2783] = 33'd3864863391;
        test_addr[2784] = 338;
        test_data[2784] = 33'd78882875;
        test_addr[2785] = 339;
        test_data[2785] = 33'd214478531;
        test_addr[2786] = 340;
        test_data[2786] = 33'd3336040161;
        test_addr[2787] = 341;
        test_data[2787] = 33'd742447467;
        test_addr[2788] = 342;
        test_data[2788] = 33'd1626249509;
        test_addr[2789] = 343;
        test_data[2789] = 33'd5532774551;
        test_addr[2790] = 344;
        test_data[2790] = 33'd281373290;
        test_addr[2791] = 345;
        test_data[2791] = 33'd3040204748;
        test_addr[2792] = 346;
        test_data[2792] = 33'd571024672;
        test_addr[2793] = 347;
        test_data[2793] = 33'd5022506074;
        test_addr[2794] = 348;
        test_data[2794] = 33'd6062446500;
        test_addr[2795] = 349;
        test_data[2795] = 33'd516820221;
        test_addr[2796] = 350;
        test_data[2796] = 33'd6262592210;
        test_addr[2797] = 351;
        test_data[2797] = 33'd1077652121;
        test_addr[2798] = 352;
        test_data[2798] = 33'd147931898;
        test_addr[2799] = 353;
        test_data[2799] = 33'd1549263986;
        test_addr[2800] = 354;
        test_data[2800] = 33'd3966319412;
        test_addr[2801] = 355;
        test_data[2801] = 33'd8542565854;
        test_addr[2802] = 356;
        test_data[2802] = 33'd7445234518;
        test_addr[2803] = 357;
        test_data[2803] = 33'd7520835263;
        test_addr[2804] = 719;
        test_data[2804] = 33'd8268833177;
        test_addr[2805] = 720;
        test_data[2805] = 33'd2104937406;
        test_addr[2806] = 721;
        test_data[2806] = 33'd1128753372;
        test_addr[2807] = 722;
        test_data[2807] = 33'd2657954045;
        test_addr[2808] = 723;
        test_data[2808] = 33'd3748128516;
        test_addr[2809] = 724;
        test_data[2809] = 33'd7936337354;
        test_addr[2810] = 725;
        test_data[2810] = 33'd1658946223;
        test_addr[2811] = 726;
        test_data[2811] = 33'd2309348786;
        test_addr[2812] = 727;
        test_data[2812] = 33'd3471679949;
        test_addr[2813] = 728;
        test_data[2813] = 33'd8059006419;
        test_addr[2814] = 729;
        test_data[2814] = 33'd919345546;
        test_addr[2815] = 730;
        test_data[2815] = 33'd4067928788;
        test_addr[2816] = 731;
        test_data[2816] = 33'd7805200090;
        test_addr[2817] = 732;
        test_data[2817] = 33'd8396419921;
        test_addr[2818] = 733;
        test_data[2818] = 33'd6730312318;
        test_addr[2819] = 734;
        test_data[2819] = 33'd7012996499;
        test_addr[2820] = 735;
        test_data[2820] = 33'd1970925193;
        test_addr[2821] = 736;
        test_data[2821] = 33'd2719855705;
        test_addr[2822] = 737;
        test_data[2822] = 33'd3147194239;
        test_addr[2823] = 738;
        test_data[2823] = 33'd4401607318;
        test_addr[2824] = 739;
        test_data[2824] = 33'd3426545964;
        test_addr[2825] = 740;
        test_data[2825] = 33'd3233147737;
        test_addr[2826] = 741;
        test_data[2826] = 33'd6629303403;
        test_addr[2827] = 742;
        test_data[2827] = 33'd4364296600;
        test_addr[2828] = 743;
        test_data[2828] = 33'd911610565;
        test_addr[2829] = 744;
        test_data[2829] = 33'd3214813081;
        test_addr[2830] = 745;
        test_data[2830] = 33'd6149777987;
        test_addr[2831] = 746;
        test_data[2831] = 33'd1275703116;
        test_addr[2832] = 358;
        test_data[2832] = 33'd928067253;
        test_addr[2833] = 359;
        test_data[2833] = 33'd4082684122;
        test_addr[2834] = 360;
        test_data[2834] = 33'd1677042253;
        test_addr[2835] = 361;
        test_data[2835] = 33'd851421913;
        test_addr[2836] = 362;
        test_data[2836] = 33'd739869624;
        test_addr[2837] = 363;
        test_data[2837] = 33'd3444286968;
        test_addr[2838] = 364;
        test_data[2838] = 33'd5354630784;
        test_addr[2839] = 365;
        test_data[2839] = 33'd1008210114;
        test_addr[2840] = 366;
        test_data[2840] = 33'd6659480754;
        test_addr[2841] = 367;
        test_data[2841] = 33'd916394114;
        test_addr[2842] = 368;
        test_data[2842] = 33'd1550869304;
        test_addr[2843] = 369;
        test_data[2843] = 33'd5020644837;
        test_addr[2844] = 370;
        test_data[2844] = 33'd4039069504;
        test_addr[2845] = 371;
        test_data[2845] = 33'd1796770481;
        test_addr[2846] = 372;
        test_data[2846] = 33'd7150280742;
        test_addr[2847] = 373;
        test_data[2847] = 33'd6943526;
        test_addr[2848] = 374;
        test_data[2848] = 33'd8299256744;
        test_addr[2849] = 375;
        test_data[2849] = 33'd6973810512;
        test_addr[2850] = 376;
        test_data[2850] = 33'd3383574487;
        test_addr[2851] = 377;
        test_data[2851] = 33'd258678087;
        test_addr[2852] = 378;
        test_data[2852] = 33'd1707274193;
        test_addr[2853] = 379;
        test_data[2853] = 33'd76696075;
        test_addr[2854] = 380;
        test_data[2854] = 33'd4157069748;
        test_addr[2855] = 381;
        test_data[2855] = 33'd3760007301;
        test_addr[2856] = 382;
        test_data[2856] = 33'd4735221545;
        test_addr[2857] = 383;
        test_data[2857] = 33'd7116307232;
        test_addr[2858] = 384;
        test_data[2858] = 33'd3879200274;
        test_addr[2859] = 385;
        test_data[2859] = 33'd1458835581;
        test_addr[2860] = 386;
        test_data[2860] = 33'd1621402957;
        test_addr[2861] = 387;
        test_data[2861] = 33'd7651392653;
        test_addr[2862] = 388;
        test_data[2862] = 33'd4716586721;
        test_addr[2863] = 389;
        test_data[2863] = 33'd691041695;
        test_addr[2864] = 390;
        test_data[2864] = 33'd5415202904;
        test_addr[2865] = 391;
        test_data[2865] = 33'd4156755592;
        test_addr[2866] = 392;
        test_data[2866] = 33'd3669726690;
        test_addr[2867] = 393;
        test_data[2867] = 33'd3584816215;
        test_addr[2868] = 394;
        test_data[2868] = 33'd5103112722;
        test_addr[2869] = 395;
        test_data[2869] = 33'd3549743356;
        test_addr[2870] = 396;
        test_data[2870] = 33'd179786261;
        test_addr[2871] = 397;
        test_data[2871] = 33'd3874668741;
        test_addr[2872] = 398;
        test_data[2872] = 33'd2124586123;
        test_addr[2873] = 399;
        test_data[2873] = 33'd8165423036;
        test_addr[2874] = 400;
        test_data[2874] = 33'd2260948046;
        test_addr[2875] = 401;
        test_data[2875] = 33'd977523721;
        test_addr[2876] = 402;
        test_data[2876] = 33'd8087271904;
        test_addr[2877] = 403;
        test_data[2877] = 33'd603897780;
        test_addr[2878] = 404;
        test_data[2878] = 33'd284306586;
        test_addr[2879] = 405;
        test_data[2879] = 33'd8213729496;
        test_addr[2880] = 406;
        test_data[2880] = 33'd8194325843;
        test_addr[2881] = 407;
        test_data[2881] = 33'd3309369165;
        test_addr[2882] = 408;
        test_data[2882] = 33'd6887144926;
        test_addr[2883] = 409;
        test_data[2883] = 33'd1708234285;
        test_addr[2884] = 410;
        test_data[2884] = 33'd5920019766;
        test_addr[2885] = 411;
        test_data[2885] = 33'd3626126882;
        test_addr[2886] = 412;
        test_data[2886] = 33'd1506882181;
        test_addr[2887] = 413;
        test_data[2887] = 33'd2482816989;
        test_addr[2888] = 414;
        test_data[2888] = 33'd7458676951;
        test_addr[2889] = 415;
        test_data[2889] = 33'd2824809495;
        test_addr[2890] = 176;
        test_data[2890] = 33'd2422858599;
        test_addr[2891] = 177;
        test_data[2891] = 33'd4706719510;
        test_addr[2892] = 178;
        test_data[2892] = 33'd745299376;
        test_addr[2893] = 179;
        test_data[2893] = 33'd7845033967;
        test_addr[2894] = 180;
        test_data[2894] = 33'd4240384840;
        test_addr[2895] = 181;
        test_data[2895] = 33'd2156248305;
        test_addr[2896] = 182;
        test_data[2896] = 33'd1222529405;
        test_addr[2897] = 416;
        test_data[2897] = 33'd2818957874;
        test_addr[2898] = 355;
        test_data[2898] = 33'd4247598558;
        test_addr[2899] = 356;
        test_data[2899] = 33'd4343062119;
        test_addr[2900] = 357;
        test_data[2900] = 33'd3225867967;
        test_addr[2901] = 358;
        test_data[2901] = 33'd928067253;
        test_addr[2902] = 359;
        test_data[2902] = 33'd4082684122;
        test_addr[2903] = 360;
        test_data[2903] = 33'd6101445514;
        test_addr[2904] = 361;
        test_data[2904] = 33'd6469415934;
        test_addr[2905] = 362;
        test_data[2905] = 33'd739869624;
        test_addr[2906] = 363;
        test_data[2906] = 33'd3444286968;
        test_addr[2907] = 364;
        test_data[2907] = 33'd8530555955;
        test_addr[2908] = 417;
        test_data[2908] = 33'd4549617601;
        test_addr[2909] = 418;
        test_data[2909] = 33'd1591263160;
        test_addr[2910] = 419;
        test_data[2910] = 33'd188335908;
        test_addr[2911] = 420;
        test_data[2911] = 33'd1107395673;
        test_addr[2912] = 421;
        test_data[2912] = 33'd4979502503;
        test_addr[2913] = 422;
        test_data[2913] = 33'd7323289186;
        test_addr[2914] = 423;
        test_data[2914] = 33'd6531454784;
        test_addr[2915] = 424;
        test_data[2915] = 33'd458707520;
        test_addr[2916] = 425;
        test_data[2916] = 33'd2344341674;
        test_addr[2917] = 426;
        test_data[2917] = 33'd1116232863;
        test_addr[2918] = 427;
        test_data[2918] = 33'd5138412184;
        test_addr[2919] = 428;
        test_data[2919] = 33'd6289407438;
        test_addr[2920] = 429;
        test_data[2920] = 33'd8016443797;
        test_addr[2921] = 430;
        test_data[2921] = 33'd4903856201;
        test_addr[2922] = 431;
        test_data[2922] = 33'd894319900;
        test_addr[2923] = 432;
        test_data[2923] = 33'd8001618907;
        test_addr[2924] = 433;
        test_data[2924] = 33'd2905210644;
        test_addr[2925] = 434;
        test_data[2925] = 33'd8490840848;
        test_addr[2926] = 435;
        test_data[2926] = 33'd1781223650;
        test_addr[2927] = 436;
        test_data[2927] = 33'd1024435444;
        test_addr[2928] = 437;
        test_data[2928] = 33'd7583645711;
        test_addr[2929] = 438;
        test_data[2929] = 33'd3957892093;
        test_addr[2930] = 439;
        test_data[2930] = 33'd5354734070;
        test_addr[2931] = 440;
        test_data[2931] = 33'd7635881620;
        test_addr[2932] = 441;
        test_data[2932] = 33'd6389302668;
        test_addr[2933] = 442;
        test_data[2933] = 33'd435473850;
        test_addr[2934] = 443;
        test_data[2934] = 33'd2309805798;
        test_addr[2935] = 444;
        test_data[2935] = 33'd239030141;
        test_addr[2936] = 445;
        test_data[2936] = 33'd57979874;
        test_addr[2937] = 446;
        test_data[2937] = 33'd185249361;
        test_addr[2938] = 447;
        test_data[2938] = 33'd6706183398;
        test_addr[2939] = 448;
        test_data[2939] = 33'd229452757;
        test_addr[2940] = 449;
        test_data[2940] = 33'd2000661367;
        test_addr[2941] = 450;
        test_data[2941] = 33'd1220832376;
        test_addr[2942] = 451;
        test_data[2942] = 33'd4533972187;
        test_addr[2943] = 452;
        test_data[2943] = 33'd6707236459;
        test_addr[2944] = 453;
        test_data[2944] = 33'd2615425596;
        test_addr[2945] = 954;
        test_data[2945] = 33'd2796648127;
        test_addr[2946] = 955;
        test_data[2946] = 33'd6158771864;
        test_addr[2947] = 956;
        test_data[2947] = 33'd90020364;
        test_addr[2948] = 957;
        test_data[2948] = 33'd2991872276;
        test_addr[2949] = 958;
        test_data[2949] = 33'd3447221745;
        test_addr[2950] = 959;
        test_data[2950] = 33'd3794599805;
        test_addr[2951] = 960;
        test_data[2951] = 33'd8198675403;
        test_addr[2952] = 454;
        test_data[2952] = 33'd2272728078;
        test_addr[2953] = 941;
        test_data[2953] = 33'd1460688612;
        test_addr[2954] = 942;
        test_data[2954] = 33'd3185997769;
        test_addr[2955] = 943;
        test_data[2955] = 33'd6551889632;
        test_addr[2956] = 944;
        test_data[2956] = 33'd1934668787;
        test_addr[2957] = 945;
        test_data[2957] = 33'd1342625013;
        test_addr[2958] = 946;
        test_data[2958] = 33'd1984305920;
        test_addr[2959] = 947;
        test_data[2959] = 33'd3397671939;
        test_addr[2960] = 948;
        test_data[2960] = 33'd689974145;
        test_addr[2961] = 949;
        test_data[2961] = 33'd5480768056;
        test_addr[2962] = 950;
        test_data[2962] = 33'd4403735772;
        test_addr[2963] = 951;
        test_data[2963] = 33'd7453723562;
        test_addr[2964] = 455;
        test_data[2964] = 33'd3050926603;
        test_addr[2965] = 296;
        test_data[2965] = 33'd4844554616;
        test_addr[2966] = 297;
        test_data[2966] = 33'd6858094358;
        test_addr[2967] = 298;
        test_data[2967] = 33'd8141418113;
        test_addr[2968] = 299;
        test_data[2968] = 33'd2163199348;
        test_addr[2969] = 300;
        test_data[2969] = 33'd1880021582;
        test_addr[2970] = 301;
        test_data[2970] = 33'd5849546378;
        test_addr[2971] = 302;
        test_data[2971] = 33'd6411323653;
        test_addr[2972] = 303;
        test_data[2972] = 33'd6369342743;
        test_addr[2973] = 304;
        test_data[2973] = 33'd460827716;
        test_addr[2974] = 305;
        test_data[2974] = 33'd1866235150;
        test_addr[2975] = 306;
        test_data[2975] = 33'd7828249656;
        test_addr[2976] = 307;
        test_data[2976] = 33'd6073380677;
        test_addr[2977] = 308;
        test_data[2977] = 33'd2611705428;
        test_addr[2978] = 456;
        test_data[2978] = 33'd1297742875;
        test_addr[2979] = 457;
        test_data[2979] = 33'd2700525639;
        test_addr[2980] = 458;
        test_data[2980] = 33'd2696971372;
        test_addr[2981] = 459;
        test_data[2981] = 33'd582707416;
        test_addr[2982] = 460;
        test_data[2982] = 33'd5323803017;
        test_addr[2983] = 461;
        test_data[2983] = 33'd583606136;
        test_addr[2984] = 462;
        test_data[2984] = 33'd3772793346;
        test_addr[2985] = 463;
        test_data[2985] = 33'd5098386797;
        test_addr[2986] = 464;
        test_data[2986] = 33'd6312812802;
        test_addr[2987] = 465;
        test_data[2987] = 33'd6715642686;
        test_addr[2988] = 466;
        test_data[2988] = 33'd2807963646;
        test_addr[2989] = 426;
        test_data[2989] = 33'd5311441109;
        test_addr[2990] = 427;
        test_data[2990] = 33'd6955347948;
        test_addr[2991] = 428;
        test_data[2991] = 33'd1994440142;
        test_addr[2992] = 429;
        test_data[2992] = 33'd3721476501;
        test_addr[2993] = 430;
        test_data[2993] = 33'd608888905;
        test_addr[2994] = 431;
        test_data[2994] = 33'd894319900;
        test_addr[2995] = 432;
        test_data[2995] = 33'd3706651611;
        test_addr[2996] = 467;
        test_data[2996] = 33'd7291179223;
        test_addr[2997] = 468;
        test_data[2997] = 33'd2873278775;
        test_addr[2998] = 469;
        test_data[2998] = 33'd4108189927;
        test_addr[2999] = 470;
        test_data[2999] = 33'd1183712898;

    end
endmodule

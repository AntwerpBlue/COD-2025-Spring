
`timescale 1ns/1ps
module mem_bram #(
    parameter ADDR_WIDTH = 10,		//地址宽度
    parameter DATA_WIDTH = 128		//数据宽度
)(
    input                   clk,   // Clock
    input [ADDR_WIDTH-1:0]  raddr,  // Address
    input [ADDR_WIDTH-1:0]  waddr,  // Address
    input [DATA_WIDTH-1:0]  din,   // Data Input
    input                   we,    // Write Enable
    output [DATA_WIDTH-1:0] dout   // Data Output
); 
    reg [ADDR_WIDTH-1:0] addr_r;  // Address Register
    reg [DATA_WIDTH-1:0] ram [0:(1 << ADDR_WIDTH)-1];
    integer i;
    initial begin
        ram[0][31:0] = 32'd2266818756;
        ram[0][63:32] = 32'd2545176946;
        ram[0][95:64] = 32'd3771999802;
        ram[0][127:96] = 32'd24445434;
        ram[1][31:0] = 32'd2235130613;
        ram[1][63:32] = 32'd2372128561;
        ram[1][95:64] = 32'd1280683540;
        ram[1][127:96] = 32'd881802803;
        ram[2][31:0] = 32'd3524160583;
        ram[2][63:32] = 32'd2731114248;
        ram[2][95:64] = 32'd3358287115;
        ram[2][127:96] = 32'd3681162206;
        ram[3][31:0] = 32'd4028186270;
        ram[3][63:32] = 32'd1541123444;
        ram[3][95:64] = 32'd1979349311;
        ram[3][127:96] = 32'd3336181142;
        ram[4][31:0] = 32'd4425813;
        ram[4][63:32] = 32'd2023586953;
        ram[4][95:64] = 32'd1691049431;
        ram[4][127:96] = 32'd2420327030;
        ram[5][31:0] = 32'd892044972;
        ram[5][63:32] = 32'd2561191935;
        ram[5][95:64] = 32'd9397193;
        ram[5][127:96] = 32'd2154342992;
        ram[6][31:0] = 32'd1503049;
        ram[6][63:32] = 32'd2605255280;
        ram[6][95:64] = 32'd385819564;
        ram[6][127:96] = 32'd3441740048;
        ram[7][31:0] = 32'd1087055728;
        ram[7][63:32] = 32'd1848244721;
        ram[7][95:64] = 32'd2237310583;
        ram[7][127:96] = 32'd1855015640;
        ram[8][31:0] = 32'd514700352;
        ram[8][63:32] = 32'd3931481952;
        ram[8][95:64] = 32'd2988630753;
        ram[8][127:96] = 32'd1427007413;
        ram[9][31:0] = 32'd2361056536;
        ram[9][63:32] = 32'd4017425673;
        ram[9][95:64] = 32'd2401565710;
        ram[9][127:96] = 32'd3097257097;
        ram[10][31:0] = 32'd2224301287;
        ram[10][63:32] = 32'd190445736;
        ram[10][95:64] = 32'd3652372969;
        ram[10][127:96] = 32'd2636643983;
        ram[11][31:0] = 32'd1301135708;
        ram[11][63:32] = 32'd2614948748;
        ram[11][95:64] = 32'd1936612333;
        ram[11][127:96] = 32'd2919107533;
        ram[12][31:0] = 32'd2774778100;
        ram[12][63:32] = 32'd751512591;
        ram[12][95:64] = 32'd3387573992;
        ram[12][127:96] = 32'd1434736929;
        ram[13][31:0] = 32'd1963808414;
        ram[13][63:32] = 32'd3378935871;
        ram[13][95:64] = 32'd2589183808;
        ram[13][127:96] = 32'd1382426006;
        ram[14][31:0] = 32'd3847507083;
        ram[14][63:32] = 32'd2855835886;
        ram[14][95:64] = 32'd2866622380;
        ram[14][127:96] = 32'd2199430969;
        ram[15][31:0] = 32'd305410629;
        ram[15][63:32] = 32'd3243858099;
        ram[15][95:64] = 32'd4196019249;
        ram[15][127:96] = 32'd100769450;
        ram[16][31:0] = 32'd3038722049;
        ram[16][63:32] = 32'd993562414;
        ram[16][95:64] = 32'd2051708468;
        ram[16][127:96] = 32'd3639768664;
        ram[17][31:0] = 32'd2031775880;
        ram[17][63:32] = 32'd1753936223;
        ram[17][95:64] = 32'd1368704711;
        ram[17][127:96] = 32'd3950328245;
        ram[18][31:0] = 32'd2563905635;
        ram[18][63:32] = 32'd220268032;
        ram[18][95:64] = 32'd3405503829;
        ram[18][127:96] = 32'd2274537304;
        ram[19][31:0] = 32'd2531899576;
        ram[19][63:32] = 32'd1279103495;
        ram[19][95:64] = 32'd258451118;
        ram[19][127:96] = 32'd3379420619;
        ram[20][31:0] = 32'd818068638;
        ram[20][63:32] = 32'd1332563736;
        ram[20][95:64] = 32'd1240469410;
        ram[20][127:96] = 32'd681728304;
        ram[21][31:0] = 32'd1553318842;
        ram[21][63:32] = 32'd3303270017;
        ram[21][95:64] = 32'd740045131;
        ram[21][127:96] = 32'd2854372909;
        ram[22][31:0] = 32'd4094716213;
        ram[22][63:32] = 32'd3855383794;
        ram[22][95:64] = 32'd4119473539;
        ram[22][127:96] = 32'd3196504029;
        ram[23][31:0] = 32'd4229662223;
        ram[23][63:32] = 32'd263550839;
        ram[23][95:64] = 32'd2300279539;
        ram[23][127:96] = 32'd2832430349;
        ram[24][31:0] = 32'd1856102477;
        ram[24][63:32] = 32'd2839264634;
        ram[24][95:64] = 32'd4210654701;
        ram[24][127:96] = 32'd2883454270;
        ram[25][31:0] = 32'd3239304748;
        ram[25][63:32] = 32'd2986556686;
        ram[25][95:64] = 32'd1124317209;
        ram[25][127:96] = 32'd2627891325;
        ram[26][31:0] = 32'd3714367826;
        ram[26][63:32] = 32'd3407001355;
        ram[26][95:64] = 32'd898134430;
        ram[26][127:96] = 32'd4243198286;
        ram[27][31:0] = 32'd52659899;
        ram[27][63:32] = 32'd2394762171;
        ram[27][95:64] = 32'd2924822209;
        ram[27][127:96] = 32'd3939766389;
        ram[28][31:0] = 32'd241897106;
        ram[28][63:32] = 32'd2590394246;
        ram[28][95:64] = 32'd3614315923;
        ram[28][127:96] = 32'd2347364473;
        ram[29][31:0] = 32'd126332533;
        ram[29][63:32] = 32'd3765837093;
        ram[29][95:64] = 32'd4130850739;
        ram[29][127:96] = 32'd1052542082;
        ram[30][31:0] = 32'd3448262298;
        ram[30][63:32] = 32'd157354656;
        ram[30][95:64] = 32'd1522076612;
        ram[30][127:96] = 32'd3515538989;
        ram[31][31:0] = 32'd563225304;
        ram[31][63:32] = 32'd2709632180;
        ram[31][95:64] = 32'd2525024090;
        ram[31][127:96] = 32'd3999854979;
        ram[32][31:0] = 32'd1320669106;
        ram[32][63:32] = 32'd4160678548;
        ram[32][95:64] = 32'd1268433295;
        ram[32][127:96] = 32'd917885500;
        ram[33][31:0] = 32'd3529417599;
        ram[33][63:32] = 32'd1645346336;
        ram[33][95:64] = 32'd2206256073;
        ram[33][127:96] = 32'd2550195621;
        ram[34][31:0] = 32'd3884710849;
        ram[34][63:32] = 32'd1980778037;
        ram[34][95:64] = 32'd2910298998;
        ram[34][127:96] = 32'd3677407724;
        ram[35][31:0] = 32'd3005608887;
        ram[35][63:32] = 32'd324907900;
        ram[35][95:64] = 32'd2983160463;
        ram[35][127:96] = 32'd796190208;
        ram[36][31:0] = 32'd4214779887;
        ram[36][63:32] = 32'd1207656834;
        ram[36][95:64] = 32'd2005652566;
        ram[36][127:96] = 32'd2764225137;
        ram[37][31:0] = 32'd3002299453;
        ram[37][63:32] = 32'd2268132089;
        ram[37][95:64] = 32'd1321807965;
        ram[37][127:96] = 32'd199031358;
        ram[38][31:0] = 32'd4105911548;
        ram[38][63:32] = 32'd632865373;
        ram[38][95:64] = 32'd1881539630;
        ram[38][127:96] = 32'd1302683176;
        ram[39][31:0] = 32'd3852022963;
        ram[39][63:32] = 32'd287346741;
        ram[39][95:64] = 32'd217812934;
        ram[39][127:96] = 32'd234338877;
        ram[40][31:0] = 32'd1681817037;
        ram[40][63:32] = 32'd914326549;
        ram[40][95:64] = 32'd1711500696;
        ram[40][127:96] = 32'd2753348300;
        ram[41][31:0] = 32'd2463360826;
        ram[41][63:32] = 32'd106644142;
        ram[41][95:64] = 32'd1831422667;
        ram[41][127:96] = 32'd188544578;
        ram[42][31:0] = 32'd547216839;
        ram[42][63:32] = 32'd1498396855;
        ram[42][95:64] = 32'd2103127943;
        ram[42][127:96] = 32'd1241383773;
        ram[43][31:0] = 32'd1555194164;
        ram[43][63:32] = 32'd1456155483;
        ram[43][95:64] = 32'd3331308539;
        ram[43][127:96] = 32'd2297598737;
        ram[44][31:0] = 32'd2275341057;
        ram[44][63:32] = 32'd2198187797;
        ram[44][95:64] = 32'd3283596447;
        ram[44][127:96] = 32'd2011666985;
        ram[45][31:0] = 32'd4026446541;
        ram[45][63:32] = 32'd2341176196;
        ram[45][95:64] = 32'd2294431329;
        ram[45][127:96] = 32'd563757395;
        ram[46][31:0] = 32'd1125354659;
        ram[46][63:32] = 32'd1560025071;
        ram[46][95:64] = 32'd3682629875;
        ram[46][127:96] = 32'd3384354663;
        ram[47][31:0] = 32'd4083814239;
        ram[47][63:32] = 32'd3994613051;
        ram[47][95:64] = 32'd2487141371;
        ram[47][127:96] = 32'd1599404350;
        ram[48][31:0] = 32'd2694434016;
        ram[48][63:32] = 32'd3086054301;
        ram[48][95:64] = 32'd2912051046;
        ram[48][127:96] = 32'd3059700818;
        ram[49][31:0] = 32'd2957372585;
        ram[49][63:32] = 32'd3763869217;
        ram[49][95:64] = 32'd4018594710;
        ram[49][127:96] = 32'd1897789635;
        ram[50][31:0] = 32'd4007449550;
        ram[50][63:32] = 32'd29735866;
        ram[50][95:64] = 32'd878548522;
        ram[50][127:96] = 32'd4132021586;
        ram[51][31:0] = 32'd3794704459;
        ram[51][63:32] = 32'd2173752367;
        ram[51][95:64] = 32'd380753888;
        ram[51][127:96] = 32'd843754471;
        ram[52][31:0] = 32'd3209549992;
        ram[52][63:32] = 32'd87559006;
        ram[52][95:64] = 32'd2782581352;
        ram[52][127:96] = 32'd3322545857;
        ram[53][31:0] = 32'd1617687132;
        ram[53][63:32] = 32'd2155161093;
        ram[53][95:64] = 32'd3250589043;
        ram[53][127:96] = 32'd1844038646;
        ram[54][31:0] = 32'd114160115;
        ram[54][63:32] = 32'd1912963371;
        ram[54][95:64] = 32'd321338277;
        ram[54][127:96] = 32'd308900539;
        ram[55][31:0] = 32'd1136133958;
        ram[55][63:32] = 32'd3414348433;
        ram[55][95:64] = 32'd1146860549;
        ram[55][127:96] = 32'd3536349469;
        ram[56][31:0] = 32'd2844672327;
        ram[56][63:32] = 32'd541535233;
        ram[56][95:64] = 32'd4004290607;
        ram[56][127:96] = 32'd905576619;
        ram[57][31:0] = 32'd3498918036;
        ram[57][63:32] = 32'd1164658069;
        ram[57][95:64] = 32'd3123327297;
        ram[57][127:96] = 32'd1147904076;
        ram[58][31:0] = 32'd930589679;
        ram[58][63:32] = 32'd1289878889;
        ram[58][95:64] = 32'd2502772052;
        ram[58][127:96] = 32'd675031687;
        ram[59][31:0] = 32'd983334167;
        ram[59][63:32] = 32'd2066899154;
        ram[59][95:64] = 32'd993254642;
        ram[59][127:96] = 32'd1377847727;
        ram[60][31:0] = 32'd3107113144;
        ram[60][63:32] = 32'd1429672039;
        ram[60][95:64] = 32'd2777853686;
        ram[60][127:96] = 32'd3048963064;
        ram[61][31:0] = 32'd1306044194;
        ram[61][63:32] = 32'd2052459312;
        ram[61][95:64] = 32'd1635138116;
        ram[61][127:96] = 32'd1963291307;
        ram[62][31:0] = 32'd810408981;
        ram[62][63:32] = 32'd3978129519;
        ram[62][95:64] = 32'd673588786;
        ram[62][127:96] = 32'd1773791810;
        ram[63][31:0] = 32'd2454902627;
        ram[63][63:32] = 32'd2796634323;
        ram[63][95:64] = 32'd4032840749;
        ram[63][127:96] = 32'd3596974217;
        ram[64][31:0] = 32'd2781187333;
        ram[64][63:32] = 32'd894384987;
        ram[64][95:64] = 32'd3514343316;
        ram[64][127:96] = 32'd3390847646;
        ram[65][31:0] = 32'd3363163059;
        ram[65][63:32] = 32'd629678269;
        ram[65][95:64] = 32'd4191130667;
        ram[65][127:96] = 32'd2580999626;
        ram[66][31:0] = 32'd687477629;
        ram[66][63:32] = 32'd3171138656;
        ram[66][95:64] = 32'd966539116;
        ram[66][127:96] = 32'd2125390319;
        ram[67][31:0] = 32'd59643427;
        ram[67][63:32] = 32'd2017951304;
        ram[67][95:64] = 32'd2409706630;
        ram[67][127:96] = 32'd2718986291;
        ram[68][31:0] = 32'd478200901;
        ram[68][63:32] = 32'd56693191;
        ram[68][95:64] = 32'd3318236443;
        ram[68][127:96] = 32'd3432839275;
        ram[69][31:0] = 32'd629857851;
        ram[69][63:32] = 32'd764865874;
        ram[69][95:64] = 32'd3400886719;
        ram[69][127:96] = 32'd3495680488;
        ram[70][31:0] = 32'd761284035;
        ram[70][63:32] = 32'd3944389777;
        ram[70][95:64] = 32'd1686295980;
        ram[70][127:96] = 32'd2681193817;
        ram[71][31:0] = 32'd2666681427;
        ram[71][63:32] = 32'd1435481041;
        ram[71][95:64] = 32'd2360048588;
        ram[71][127:96] = 32'd3189797644;
        ram[72][31:0] = 32'd2754042220;
        ram[72][63:32] = 32'd3204524255;
        ram[72][95:64] = 32'd3989670362;
        ram[72][127:96] = 32'd3655503747;
        ram[73][31:0] = 32'd2039041372;
        ram[73][63:32] = 32'd3750343722;
        ram[73][95:64] = 32'd228860212;
        ram[73][127:96] = 32'd811886581;
        ram[74][31:0] = 32'd262993620;
        ram[74][63:32] = 32'd2277946841;
        ram[74][95:64] = 32'd1530159267;
        ram[74][127:96] = 32'd3707209855;
        ram[75][31:0] = 32'd2615739423;
        ram[75][63:32] = 32'd3075188539;
        ram[75][95:64] = 32'd35142408;
        ram[75][127:96] = 32'd143048814;
        ram[76][31:0] = 32'd3014575534;
        ram[76][63:32] = 32'd2393483621;
        ram[76][95:64] = 32'd1818292495;
        ram[76][127:96] = 32'd2982069157;
        ram[77][31:0] = 32'd2458562695;
        ram[77][63:32] = 32'd714351707;
        ram[77][95:64] = 32'd3692301779;
        ram[77][127:96] = 32'd3880279301;
        ram[78][31:0] = 32'd1985873362;
        ram[78][63:32] = 32'd362309121;
        ram[78][95:64] = 32'd751501571;
        ram[78][127:96] = 32'd1263301752;
        ram[79][31:0] = 32'd3154340319;
        ram[79][63:32] = 32'd631004568;
        ram[79][95:64] = 32'd3901681998;
        ram[79][127:96] = 32'd2331515849;
        ram[80][31:0] = 32'd3248669603;
        ram[80][63:32] = 32'd2361956255;
        ram[80][95:64] = 32'd3243207308;
        ram[80][127:96] = 32'd1882614181;
        ram[81][31:0] = 32'd330852185;
        ram[81][63:32] = 32'd539824620;
        ram[81][95:64] = 32'd2972100094;
        ram[81][127:96] = 32'd1156839342;
        ram[82][31:0] = 32'd952282828;
        ram[82][63:32] = 32'd3903899561;
        ram[82][95:64] = 32'd2287195610;
        ram[82][127:96] = 32'd3237563871;
        ram[83][31:0] = 32'd2406902933;
        ram[83][63:32] = 32'd509475252;
        ram[83][95:64] = 32'd3431054307;
        ram[83][127:96] = 32'd241135054;
        ram[84][31:0] = 32'd3346235914;
        ram[84][63:32] = 32'd1691010132;
        ram[84][95:64] = 32'd3573453669;
        ram[84][127:96] = 32'd944678627;
        ram[85][31:0] = 32'd3309872861;
        ram[85][63:32] = 32'd3239124403;
        ram[85][95:64] = 32'd744650674;
        ram[85][127:96] = 32'd2055667857;
        ram[86][31:0] = 32'd253890222;
        ram[86][63:32] = 32'd2662284645;
        ram[86][95:64] = 32'd3114256567;
        ram[86][127:96] = 32'd2552236765;
        ram[87][31:0] = 32'd3765498237;
        ram[87][63:32] = 32'd2317422068;
        ram[87][95:64] = 32'd3946888309;
        ram[87][127:96] = 32'd296741918;
        ram[88][31:0] = 32'd3944142242;
        ram[88][63:32] = 32'd3399552858;
        ram[88][95:64] = 32'd2820300650;
        ram[88][127:96] = 32'd3862589515;
        ram[89][31:0] = 32'd2587005368;
        ram[89][63:32] = 32'd4022908127;
        ram[89][95:64] = 32'd3979567529;
        ram[89][127:96] = 32'd3691641483;
        ram[90][31:0] = 32'd3609013038;
        ram[90][63:32] = 32'd3669843007;
        ram[90][95:64] = 32'd4225808861;
        ram[90][127:96] = 32'd2176499912;
        ram[91][31:0] = 32'd4222053268;
        ram[91][63:32] = 32'd369210451;
        ram[91][95:64] = 32'd648433376;
        ram[91][127:96] = 32'd3620341239;
        ram[92][31:0] = 32'd3346930613;
        ram[92][63:32] = 32'd1161521471;
        ram[92][95:64] = 32'd469255750;
        ram[92][127:96] = 32'd941454407;
        ram[93][31:0] = 32'd3706783982;
        ram[93][63:32] = 32'd2520742008;
        ram[93][95:64] = 32'd2011634502;
        ram[93][127:96] = 32'd1408822660;
        ram[94][31:0] = 32'd3017136644;
        ram[94][63:32] = 32'd2966812082;
        ram[94][95:64] = 32'd2059550719;
        ram[94][127:96] = 32'd1897669063;
        ram[95][31:0] = 32'd1024754085;
        ram[95][63:32] = 32'd3910801142;
        ram[95][95:64] = 32'd3179486996;
        ram[95][127:96] = 32'd710319605;
        ram[96][31:0] = 32'd2518713733;
        ram[96][63:32] = 32'd257588625;
        ram[96][95:64] = 32'd3669660999;
        ram[96][127:96] = 32'd984172897;
        ram[97][31:0] = 32'd378350442;
        ram[97][63:32] = 32'd2549642068;
        ram[97][95:64] = 32'd909123417;
        ram[97][127:96] = 32'd2934085416;
        ram[98][31:0] = 32'd1564494824;
        ram[98][63:32] = 32'd399811056;
        ram[98][95:64] = 32'd496284610;
        ram[98][127:96] = 32'd1292390397;
        ram[99][31:0] = 32'd2322691786;
        ram[99][63:32] = 32'd2724761539;
        ram[99][95:64] = 32'd1175204693;
        ram[99][127:96] = 32'd1875700461;
        ram[100][31:0] = 32'd545504374;
        ram[100][63:32] = 32'd3417198120;
        ram[100][95:64] = 32'd1208032225;
        ram[100][127:96] = 32'd940483063;
        ram[101][31:0] = 32'd2626802031;
        ram[101][63:32] = 32'd2226632309;
        ram[101][95:64] = 32'd1667658830;
        ram[101][127:96] = 32'd1117760925;
        ram[102][31:0] = 32'd676726005;
        ram[102][63:32] = 32'd3340352858;
        ram[102][95:64] = 32'd3405405453;
        ram[102][127:96] = 32'd3762034742;
        ram[103][31:0] = 32'd3829988349;
        ram[103][63:32] = 32'd3563808226;
        ram[103][95:64] = 32'd402300966;
        ram[103][127:96] = 32'd330435490;
        ram[104][31:0] = 32'd3819993292;
        ram[104][63:32] = 32'd1438411843;
        ram[104][95:64] = 32'd564521412;
        ram[104][127:96] = 32'd4133168253;
        ram[105][31:0] = 32'd3817791626;
        ram[105][63:32] = 32'd2522318236;
        ram[105][95:64] = 32'd4144807526;
        ram[105][127:96] = 32'd2094691022;
        ram[106][31:0] = 32'd710281784;
        ram[106][63:32] = 32'd3540322948;
        ram[106][95:64] = 32'd705611193;
        ram[106][127:96] = 32'd3998550133;
        ram[107][31:0] = 32'd1801007473;
        ram[107][63:32] = 32'd3992289899;
        ram[107][95:64] = 32'd3947540049;
        ram[107][127:96] = 32'd3304810659;
        ram[108][31:0] = 32'd926426471;
        ram[108][63:32] = 32'd4013542089;
        ram[108][95:64] = 32'd188263586;
        ram[108][127:96] = 32'd3843532341;
        ram[109][31:0] = 32'd1971182400;
        ram[109][63:32] = 32'd3188866646;
        ram[109][95:64] = 32'd2860390341;
        ram[109][127:96] = 32'd1333283651;
        ram[110][31:0] = 32'd2125874662;
        ram[110][63:32] = 32'd1603229292;
        ram[110][95:64] = 32'd1682936301;
        ram[110][127:96] = 32'd170511464;
        ram[111][31:0] = 32'd2124914818;
        ram[111][63:32] = 32'd119278519;
        ram[111][95:64] = 32'd3099163608;
        ram[111][127:96] = 32'd374939133;
        ram[112][31:0] = 32'd2388061351;
        ram[112][63:32] = 32'd1443761105;
        ram[112][95:64] = 32'd2461350224;
        ram[112][127:96] = 32'd317087304;
        ram[113][31:0] = 32'd302438381;
        ram[113][63:32] = 32'd3723143858;
        ram[113][95:64] = 32'd3130965914;
        ram[113][127:96] = 32'd2867352729;
        ram[114][31:0] = 32'd3608555727;
        ram[114][63:32] = 32'd4213395215;
        ram[114][95:64] = 32'd3114864730;
        ram[114][127:96] = 32'd2890618210;
        ram[115][31:0] = 32'd685908480;
        ram[115][63:32] = 32'd232425237;
        ram[115][95:64] = 32'd3368580872;
        ram[115][127:96] = 32'd1603013143;
        ram[116][31:0] = 32'd1561543919;
        ram[116][63:32] = 32'd2880986098;
        ram[116][95:64] = 32'd633115602;
        ram[116][127:96] = 32'd533773563;
        ram[117][31:0] = 32'd2002255513;
        ram[117][63:32] = 32'd479190319;
        ram[117][95:64] = 32'd3794027735;
        ram[117][127:96] = 32'd1336088425;
        ram[118][31:0] = 32'd2925733218;
        ram[118][63:32] = 32'd3843447121;
        ram[118][95:64] = 32'd4127845043;
        ram[118][127:96] = 32'd2883836476;
        ram[119][31:0] = 32'd3010424531;
        ram[119][63:32] = 32'd2823642870;
        ram[119][95:64] = 32'd1090530905;
        ram[119][127:96] = 32'd3763673002;
        ram[120][31:0] = 32'd648309832;
        ram[120][63:32] = 32'd3166725598;
        ram[120][95:64] = 32'd1173410456;
        ram[120][127:96] = 32'd1178549137;
        ram[121][31:0] = 32'd953158137;
        ram[121][63:32] = 32'd198421201;
        ram[121][95:64] = 32'd2789818792;
        ram[121][127:96] = 32'd3574805294;
        ram[122][31:0] = 32'd2484186896;
        ram[122][63:32] = 32'd1370496534;
        ram[122][95:64] = 32'd755275238;
        ram[122][127:96] = 32'd2211071192;
        ram[123][31:0] = 32'd2984910114;
        ram[123][63:32] = 32'd392841551;
        ram[123][95:64] = 32'd1192454332;
        ram[123][127:96] = 32'd885613252;
        ram[124][31:0] = 32'd1048502686;
        ram[124][63:32] = 32'd2590240532;
        ram[124][95:64] = 32'd3649231511;
        ram[124][127:96] = 32'd4266444285;
        ram[125][31:0] = 32'd1951278430;
        ram[125][63:32] = 32'd481823011;
        ram[125][95:64] = 32'd938899533;
        ram[125][127:96] = 32'd2825090233;
        ram[126][31:0] = 32'd2373341895;
        ram[126][63:32] = 32'd891871093;
        ram[126][95:64] = 32'd644403250;
        ram[126][127:96] = 32'd3857079307;
        ram[127][31:0] = 32'd2569124247;
        ram[127][63:32] = 32'd1404134308;
        ram[127][95:64] = 32'd363583401;
        ram[127][127:96] = 32'd308446067;
        ram[128][31:0] = 32'd112430786;
        ram[128][63:32] = 32'd3149345860;
        ram[128][95:64] = 32'd1968356132;
        ram[128][127:96] = 32'd1989592525;
        ram[129][31:0] = 32'd1259652408;
        ram[129][63:32] = 32'd385111081;
        ram[129][95:64] = 32'd856602084;
        ram[129][127:96] = 32'd1283402259;
        ram[130][31:0] = 32'd3687095609;
        ram[130][63:32] = 32'd3462858656;
        ram[130][95:64] = 32'd856211726;
        ram[130][127:96] = 32'd2266066473;
        ram[131][31:0] = 32'd1899487675;
        ram[131][63:32] = 32'd2109471715;
        ram[131][95:64] = 32'd3442288853;
        ram[131][127:96] = 32'd1169423377;
        ram[132][31:0] = 32'd3121538625;
        ram[132][63:32] = 32'd441795688;
        ram[132][95:64] = 32'd1460669932;
        ram[132][127:96] = 32'd3479564107;
        ram[133][31:0] = 32'd27322558;
        ram[133][63:32] = 32'd2689141762;
        ram[133][95:64] = 32'd1059137997;
        ram[133][127:96] = 32'd1384824159;
        ram[134][31:0] = 32'd2903832397;
        ram[134][63:32] = 32'd810473933;
        ram[134][95:64] = 32'd1157057488;
        ram[134][127:96] = 32'd4282938108;
        ram[135][31:0] = 32'd432267239;
        ram[135][63:32] = 32'd3190117241;
        ram[135][95:64] = 32'd541812541;
        ram[135][127:96] = 32'd414310236;
        ram[136][31:0] = 32'd558981164;
        ram[136][63:32] = 32'd3465705991;
        ram[136][95:64] = 32'd2040323625;
        ram[136][127:96] = 32'd2109417922;
        ram[137][31:0] = 32'd2835990504;
        ram[137][63:32] = 32'd1921589746;
        ram[137][95:64] = 32'd2861464618;
        ram[137][127:96] = 32'd3506973174;
        ram[138][31:0] = 32'd1578074022;
        ram[138][63:32] = 32'd4101269385;
        ram[138][95:64] = 32'd302584709;
        ram[138][127:96] = 32'd920282072;
        ram[139][31:0] = 32'd2629206974;
        ram[139][63:32] = 32'd2738136578;
        ram[139][95:64] = 32'd3650811963;
        ram[139][127:96] = 32'd3112428785;
        ram[140][31:0] = 32'd3890402307;
        ram[140][63:32] = 32'd3925762609;
        ram[140][95:64] = 32'd2421663304;
        ram[140][127:96] = 32'd4151707470;
        ram[141][31:0] = 32'd2994986731;
        ram[141][63:32] = 32'd2785894461;
        ram[141][95:64] = 32'd770002620;
        ram[141][127:96] = 32'd806218001;
        ram[142][31:0] = 32'd2796273124;
        ram[142][63:32] = 32'd2585983587;
        ram[142][95:64] = 32'd1501919528;
        ram[142][127:96] = 32'd2429770854;
        ram[143][31:0] = 32'd2337695322;
        ram[143][63:32] = 32'd3693245975;
        ram[143][95:64] = 32'd2900017555;
        ram[143][127:96] = 32'd402074161;
        ram[144][31:0] = 32'd2373603425;
        ram[144][63:32] = 32'd2764308383;
        ram[144][95:64] = 32'd3885536651;
        ram[144][127:96] = 32'd2718604588;
        ram[145][31:0] = 32'd436662051;
        ram[145][63:32] = 32'd4026244432;
        ram[145][95:64] = 32'd3211321851;
        ram[145][127:96] = 32'd4069883337;
        ram[146][31:0] = 32'd3681182924;
        ram[146][63:32] = 32'd3586969900;
        ram[146][95:64] = 32'd3378604480;
        ram[146][127:96] = 32'd702014159;
        ram[147][31:0] = 32'd1964315406;
        ram[147][63:32] = 32'd1283209101;
        ram[147][95:64] = 32'd2472321525;
        ram[147][127:96] = 32'd4087477473;
        ram[148][31:0] = 32'd3006473031;
        ram[148][63:32] = 32'd3555664192;
        ram[148][95:64] = 32'd3790697293;
        ram[148][127:96] = 32'd1438576721;
        ram[149][31:0] = 32'd4087896024;
        ram[149][63:32] = 32'd572393240;
        ram[149][95:64] = 32'd3684002157;
        ram[149][127:96] = 32'd275103565;
        ram[150][31:0] = 32'd1402039586;
        ram[150][63:32] = 32'd2919076942;
        ram[150][95:64] = 32'd2312199791;
        ram[150][127:96] = 32'd2447831809;
        ram[151][31:0] = 32'd70723367;
        ram[151][63:32] = 32'd1980249529;
        ram[151][95:64] = 32'd4026351905;
        ram[151][127:96] = 32'd2060971912;
        ram[152][31:0] = 32'd3331304004;
        ram[152][63:32] = 32'd4261696303;
        ram[152][95:64] = 32'd2772553067;
        ram[152][127:96] = 32'd2223272245;
        ram[153][31:0] = 32'd1651535654;
        ram[153][63:32] = 32'd2948008537;
        ram[153][95:64] = 32'd58076955;
        ram[153][127:96] = 32'd2136755942;
        ram[154][31:0] = 32'd2000952156;
        ram[154][63:32] = 32'd4244853482;
        ram[154][95:64] = 32'd2216340945;
        ram[154][127:96] = 32'd1927924971;
        ram[155][31:0] = 32'd3168866381;
        ram[155][63:32] = 32'd1890719812;
        ram[155][95:64] = 32'd2596836443;
        ram[155][127:96] = 32'd2390285345;
        ram[156][31:0] = 32'd1834205843;
        ram[156][63:32] = 32'd911987830;
        ram[156][95:64] = 32'd1808868451;
        ram[156][127:96] = 32'd3885840227;
        ram[157][31:0] = 32'd765385840;
        ram[157][63:32] = 32'd1773980868;
        ram[157][95:64] = 32'd1061389955;
        ram[157][127:96] = 32'd3451386011;
        ram[158][31:0] = 32'd162213990;
        ram[158][63:32] = 32'd3083058234;
        ram[158][95:64] = 32'd2731773946;
        ram[158][127:96] = 32'd604312534;
        ram[159][31:0] = 32'd3726205383;
        ram[159][63:32] = 32'd1672692856;
        ram[159][95:64] = 32'd347823587;
        ram[159][127:96] = 32'd382292317;
        ram[160][31:0] = 32'd3936457932;
        ram[160][63:32] = 32'd1262873621;
        ram[160][95:64] = 32'd3377306771;
        ram[160][127:96] = 32'd3695691318;
        ram[161][31:0] = 32'd2891296853;
        ram[161][63:32] = 32'd543326322;
        ram[161][95:64] = 32'd1946843870;
        ram[161][127:96] = 32'd738418394;
        ram[162][31:0] = 32'd3950060224;
        ram[162][63:32] = 32'd2402313754;
        ram[162][95:64] = 32'd2885272839;
        ram[162][127:96] = 32'd1815633715;
        ram[163][31:0] = 32'd2524346705;
        ram[163][63:32] = 32'd622763873;
        ram[163][95:64] = 32'd1773452330;
        ram[163][127:96] = 32'd2678884701;
        ram[164][31:0] = 32'd2637048261;
        ram[164][63:32] = 32'd3120162192;
        ram[164][95:64] = 32'd1268986357;
        ram[164][127:96] = 32'd2764015169;
        ram[165][31:0] = 32'd3513008076;
        ram[165][63:32] = 32'd981018742;
        ram[165][95:64] = 32'd1436525592;
        ram[165][127:96] = 32'd1455377357;
        ram[166][31:0] = 32'd1694872111;
        ram[166][63:32] = 32'd1128756264;
        ram[166][95:64] = 32'd2186951376;
        ram[166][127:96] = 32'd3561967518;
        ram[167][31:0] = 32'd977172141;
        ram[167][63:32] = 32'd2603095900;
        ram[167][95:64] = 32'd2862755966;
        ram[167][127:96] = 32'd565008109;
        ram[168][31:0] = 32'd3252626599;
        ram[168][63:32] = 32'd41814705;
        ram[168][95:64] = 32'd2656360569;
        ram[168][127:96] = 32'd140747614;
        ram[169][31:0] = 32'd1174454579;
        ram[169][63:32] = 32'd4086784515;
        ram[169][95:64] = 32'd2022273082;
        ram[169][127:96] = 32'd2430705980;
        ram[170][31:0] = 32'd1235546534;
        ram[170][63:32] = 32'd1893449825;
        ram[170][95:64] = 32'd1156168669;
        ram[170][127:96] = 32'd3865309988;
        ram[171][31:0] = 32'd3058060985;
        ram[171][63:32] = 32'd4026500536;
        ram[171][95:64] = 32'd318457616;
        ram[171][127:96] = 32'd1000461927;
        ram[172][31:0] = 32'd4133517367;
        ram[172][63:32] = 32'd1681318426;
        ram[172][95:64] = 32'd4095690594;
        ram[172][127:96] = 32'd2703643781;
        ram[173][31:0] = 32'd639839837;
        ram[173][63:32] = 32'd2069998988;
        ram[173][95:64] = 32'd240080374;
        ram[173][127:96] = 32'd2186911345;
        ram[174][31:0] = 32'd2694337344;
        ram[174][63:32] = 32'd3089205481;
        ram[174][95:64] = 32'd4133583925;
        ram[174][127:96] = 32'd716758767;
        ram[175][31:0] = 32'd1777242325;
        ram[175][63:32] = 32'd1240277389;
        ram[175][95:64] = 32'd3866435097;
        ram[175][127:96] = 32'd45914204;
        ram[176][31:0] = 32'd2320769301;
        ram[176][63:32] = 32'd1506519041;
        ram[176][95:64] = 32'd2717964375;
        ram[176][127:96] = 32'd982366389;
        ram[177][31:0] = 32'd3569800214;
        ram[177][63:32] = 32'd1267071129;
        ram[177][95:64] = 32'd1657230945;
        ram[177][127:96] = 32'd2297538283;
        ram[178][31:0] = 32'd1104352139;
        ram[178][63:32] = 32'd333588719;
        ram[178][95:64] = 32'd761390289;
        ram[178][127:96] = 32'd3660057142;
        ram[179][31:0] = 32'd2391069686;
        ram[179][63:32] = 32'd2912310291;
        ram[179][95:64] = 32'd2587264415;
        ram[179][127:96] = 32'd2763934168;
        ram[180][31:0] = 32'd2954885626;
        ram[180][63:32] = 32'd1816200205;
        ram[180][95:64] = 32'd4149935825;
        ram[180][127:96] = 32'd3774650290;
        ram[181][31:0] = 32'd2475940892;
        ram[181][63:32] = 32'd711144041;
        ram[181][95:64] = 32'd3735077429;
        ram[181][127:96] = 32'd2717525231;
        ram[182][31:0] = 32'd128590783;
        ram[182][63:32] = 32'd1035742076;
        ram[182][95:64] = 32'd2774040910;
        ram[182][127:96] = 32'd1134545885;
        ram[183][31:0] = 32'd3346690204;
        ram[183][63:32] = 32'd3630483947;
        ram[183][95:64] = 32'd3464739256;
        ram[183][127:96] = 32'd2273990042;
        ram[184][31:0] = 32'd65646729;
        ram[184][63:32] = 32'd3825165600;
        ram[184][95:64] = 32'd1085936134;
        ram[184][127:96] = 32'd3116617757;
        ram[185][31:0] = 32'd2129383015;
        ram[185][63:32] = 32'd3239258243;
        ram[185][95:64] = 32'd2915364435;
        ram[185][127:96] = 32'd4186400981;
        ram[186][31:0] = 32'd912759237;
        ram[186][63:32] = 32'd469000044;
        ram[186][95:64] = 32'd2332255621;
        ram[186][127:96] = 32'd1985407323;
        ram[187][31:0] = 32'd803782110;
        ram[187][63:32] = 32'd726857318;
        ram[187][95:64] = 32'd788676881;
        ram[187][127:96] = 32'd928863370;
        ram[188][31:0] = 32'd811875741;
        ram[188][63:32] = 32'd2680759815;
        ram[188][95:64] = 32'd1886588615;
        ram[188][127:96] = 32'd2070820228;
        ram[189][31:0] = 32'd474173468;
        ram[189][63:32] = 32'd3331735711;
        ram[189][95:64] = 32'd879054465;
        ram[189][127:96] = 32'd3971751873;
        ram[190][31:0] = 32'd4199067864;
        ram[190][63:32] = 32'd2774007604;
        ram[190][95:64] = 32'd2121417843;
        ram[190][127:96] = 32'd2244486544;
        ram[191][31:0] = 32'd3976880208;
        ram[191][63:32] = 32'd1407724005;
        ram[191][95:64] = 32'd1605852982;
        ram[191][127:96] = 32'd2856339055;
        ram[192][31:0] = 32'd3795726059;
        ram[192][63:32] = 32'd3813893202;
        ram[192][95:64] = 32'd2235392260;
        ram[192][127:96] = 32'd1051449033;
        ram[193][31:0] = 32'd3678900751;
        ram[193][63:32] = 32'd2884864817;
        ram[193][95:64] = 32'd197646308;
        ram[193][127:96] = 32'd1850350391;
        ram[194][31:0] = 32'd769284591;
        ram[194][63:32] = 32'd485989889;
        ram[194][95:64] = 32'd3444963042;
        ram[194][127:96] = 32'd2260017456;
        ram[195][31:0] = 32'd404411201;
        ram[195][63:32] = 32'd2061765198;
        ram[195][95:64] = 32'd2130717397;
        ram[195][127:96] = 32'd2573492496;
        ram[196][31:0] = 32'd4161914853;
        ram[196][63:32] = 32'd1401173062;
        ram[196][95:64] = 32'd2790845645;
        ram[196][127:96] = 32'd1935616810;
        ram[197][31:0] = 32'd3121816568;
        ram[197][63:32] = 32'd2899379877;
        ram[197][95:64] = 32'd2574731272;
        ram[197][127:96] = 32'd2834578210;
        ram[198][31:0] = 32'd4103913134;
        ram[198][63:32] = 32'd1650429696;
        ram[198][95:64] = 32'd3400461738;
        ram[198][127:96] = 32'd4067395061;
        ram[199][31:0] = 32'd4142487238;
        ram[199][63:32] = 32'd2090589244;
        ram[199][95:64] = 32'd186440542;
        ram[199][127:96] = 32'd3954575845;
        ram[200][31:0] = 32'd2470310901;
        ram[200][63:32] = 32'd2849035483;
        ram[200][95:64] = 32'd4043263593;
        ram[200][127:96] = 32'd1913165819;
        ram[201][31:0] = 32'd2469310094;
        ram[201][63:32] = 32'd692126376;
        ram[201][95:64] = 32'd2817034588;
        ram[201][127:96] = 32'd2465883927;
        ram[202][31:0] = 32'd1748355561;
        ram[202][63:32] = 32'd3761030308;
        ram[202][95:64] = 32'd1557606680;
        ram[202][127:96] = 32'd712960676;
        ram[203][31:0] = 32'd2625492882;
        ram[203][63:32] = 32'd350957292;
        ram[203][95:64] = 32'd662516995;
        ram[203][127:96] = 32'd1640602374;
        ram[204][31:0] = 32'd912381185;
        ram[204][63:32] = 32'd3157715753;
        ram[204][95:64] = 32'd2986767408;
        ram[204][127:96] = 32'd1290062431;
        ram[205][31:0] = 32'd4175331955;
        ram[205][63:32] = 32'd1331449937;
        ram[205][95:64] = 32'd534736813;
        ram[205][127:96] = 32'd1932951958;
        ram[206][31:0] = 32'd3205965066;
        ram[206][63:32] = 32'd1248929761;
        ram[206][95:64] = 32'd87152189;
        ram[206][127:96] = 32'd4136395276;
        ram[207][31:0] = 32'd3880368428;
        ram[207][63:32] = 32'd1050517140;
        ram[207][95:64] = 32'd2069122430;
        ram[207][127:96] = 32'd992727670;
        ram[208][31:0] = 32'd351971474;
        ram[208][63:32] = 32'd2243381561;
        ram[208][95:64] = 32'd2798493766;
        ram[208][127:96] = 32'd3461985819;
        ram[209][31:0] = 32'd1052769268;
        ram[209][63:32] = 32'd1102094417;
        ram[209][95:64] = 32'd1113939390;
        ram[209][127:96] = 32'd851922951;
        ram[210][31:0] = 32'd3001816220;
        ram[210][63:32] = 32'd124879403;
        ram[210][95:64] = 32'd2581989200;
        ram[210][127:96] = 32'd3960620255;
        ram[211][31:0] = 32'd1272998109;
        ram[211][63:32] = 32'd2293914385;
        ram[211][95:64] = 32'd2522284635;
        ram[211][127:96] = 32'd196428976;
        ram[212][31:0] = 32'd415536288;
        ram[212][63:32] = 32'd2512243501;
        ram[212][95:64] = 32'd640217809;
        ram[212][127:96] = 32'd550630034;
        ram[213][31:0] = 32'd2146286006;
        ram[213][63:32] = 32'd3563811643;
        ram[213][95:64] = 32'd2260897852;
        ram[213][127:96] = 32'd4260287046;
        ram[214][31:0] = 32'd975862316;
        ram[214][63:32] = 32'd2261474441;
        ram[214][95:64] = 32'd2562306931;
        ram[214][127:96] = 32'd1314706587;
        ram[215][31:0] = 32'd1612728766;
        ram[215][63:32] = 32'd1715733562;
        ram[215][95:64] = 32'd1933568123;
        ram[215][127:96] = 32'd1325550564;
        ram[216][31:0] = 32'd1571587926;
        ram[216][63:32] = 32'd1605398418;
        ram[216][95:64] = 32'd3574629408;
        ram[216][127:96] = 32'd18555133;
        ram[217][31:0] = 32'd2528507951;
        ram[217][63:32] = 32'd4289214145;
        ram[217][95:64] = 32'd2749033820;
        ram[217][127:96] = 32'd3173545540;
        ram[218][31:0] = 32'd3871519302;
        ram[218][63:32] = 32'd722926779;
        ram[218][95:64] = 32'd2931664417;
        ram[218][127:96] = 32'd1365543345;
        ram[219][31:0] = 32'd3739044357;
        ram[219][63:32] = 32'd188070949;
        ram[219][95:64] = 32'd1973087823;
        ram[219][127:96] = 32'd2227416794;
        ram[220][31:0] = 32'd1923216062;
        ram[220][63:32] = 32'd554101517;
        ram[220][95:64] = 32'd4205936978;
        ram[220][127:96] = 32'd807592621;
        ram[221][31:0] = 32'd1323552558;
        ram[221][63:32] = 32'd728215166;
        ram[221][95:64] = 32'd4267669502;
        ram[221][127:96] = 32'd488449439;
        ram[222][31:0] = 32'd1386718648;
        ram[222][63:32] = 32'd4219193718;
        ram[222][95:64] = 32'd1689472630;
        ram[222][127:96] = 32'd2148240711;
        ram[223][31:0] = 32'd1634418850;
        ram[223][63:32] = 32'd3957452986;
        ram[223][95:64] = 32'd2910906105;
        ram[223][127:96] = 32'd2540543346;
        ram[224][31:0] = 32'd1587810922;
        ram[224][63:32] = 32'd2229529488;
        ram[224][95:64] = 32'd1198258543;
        ram[224][127:96] = 32'd3868985293;
        ram[225][31:0] = 32'd4008386229;
        ram[225][63:32] = 32'd3791968021;
        ram[225][95:64] = 32'd3375074483;
        ram[225][127:96] = 32'd2634020074;
        ram[226][31:0] = 32'd580095324;
        ram[226][63:32] = 32'd3362997925;
        ram[226][95:64] = 32'd1312679890;
        ram[226][127:96] = 32'd4168846095;
        ram[227][31:0] = 32'd1044409057;
        ram[227][63:32] = 32'd2141004463;
        ram[227][95:64] = 32'd4293745703;
        ram[227][127:96] = 32'd546441557;
        ram[228][31:0] = 32'd1978461553;
        ram[228][63:32] = 32'd2312966920;
        ram[228][95:64] = 32'd3697790821;
        ram[228][127:96] = 32'd1268898235;
        ram[229][31:0] = 32'd1736915697;
        ram[229][63:32] = 32'd54434874;
        ram[229][95:64] = 32'd2681524291;
        ram[229][127:96] = 32'd103226767;
        ram[230][31:0] = 32'd3925196331;
        ram[230][63:32] = 32'd680034433;
        ram[230][95:64] = 32'd715587172;
        ram[230][127:96] = 32'd4284136508;
        ram[231][31:0] = 32'd4107550478;
        ram[231][63:32] = 32'd3849164902;
        ram[231][95:64] = 32'd940863416;
        ram[231][127:96] = 32'd1927721038;
        ram[232][31:0] = 32'd2715628160;
        ram[232][63:32] = 32'd2947338001;
        ram[232][95:64] = 32'd890973601;
        ram[232][127:96] = 32'd2803979244;
        ram[233][31:0] = 32'd1290708529;
        ram[233][63:32] = 32'd2246106299;
        ram[233][95:64] = 32'd2539789535;
        ram[233][127:96] = 32'd3780989929;
        ram[234][31:0] = 32'd93762480;
        ram[234][63:32] = 32'd3186542920;
        ram[234][95:64] = 32'd1132511786;
        ram[234][127:96] = 32'd536731119;
        ram[235][31:0] = 32'd2787861430;
        ram[235][63:32] = 32'd3244851306;
        ram[235][95:64] = 32'd3431047556;
        ram[235][127:96] = 32'd1562112129;
        ram[236][31:0] = 32'd3282884071;
        ram[236][63:32] = 32'd1668354931;
        ram[236][95:64] = 32'd2538911408;
        ram[236][127:96] = 32'd965247601;
        ram[237][31:0] = 32'd4048222437;
        ram[237][63:32] = 32'd1458535013;
        ram[237][95:64] = 32'd478080935;
        ram[237][127:96] = 32'd2426414220;
        ram[238][31:0] = 32'd702855526;
        ram[238][63:32] = 32'd2168232723;
        ram[238][95:64] = 32'd2178384358;
        ram[238][127:96] = 32'd4217331207;
        ram[239][31:0] = 32'd3817405510;
        ram[239][63:32] = 32'd449348160;
        ram[239][95:64] = 32'd3257284543;
        ram[239][127:96] = 32'd3913949685;
        ram[240][31:0] = 32'd63460066;
        ram[240][63:32] = 32'd2071565022;
        ram[240][95:64] = 32'd3905065194;
        ram[240][127:96] = 32'd2423315520;
        ram[241][31:0] = 32'd1077138145;
        ram[241][63:32] = 32'd2618802793;
        ram[241][95:64] = 32'd1835137690;
        ram[241][127:96] = 32'd3880369406;
        ram[242][31:0] = 32'd3570024988;
        ram[242][63:32] = 32'd2249605407;
        ram[242][95:64] = 32'd1829669242;
        ram[242][127:96] = 32'd634864571;
        ram[243][31:0] = 32'd2410230640;
        ram[243][63:32] = 32'd2136543180;
        ram[243][95:64] = 32'd2073535736;
        ram[243][127:96] = 32'd1888922706;
        ram[244][31:0] = 32'd3839524366;
        ram[244][63:32] = 32'd1687923687;
        ram[244][95:64] = 32'd1824158172;
        ram[244][127:96] = 32'd3135075387;
        ram[245][31:0] = 32'd2435006134;
        ram[245][63:32] = 32'd250591934;
        ram[245][95:64] = 32'd772091063;
        ram[245][127:96] = 32'd509354105;
        ram[246][31:0] = 32'd1155886029;
        ram[246][63:32] = 32'd2974518957;
        ram[246][95:64] = 32'd2146402555;
        ram[246][127:96] = 32'd2638167156;
        ram[247][31:0] = 32'd3130683923;
        ram[247][63:32] = 32'd423123939;
        ram[247][95:64] = 32'd4082014275;
        ram[247][127:96] = 32'd3554038044;
        ram[248][31:0] = 32'd960033243;
        ram[248][63:32] = 32'd2909818976;
        ram[248][95:64] = 32'd1748031385;
        ram[248][127:96] = 32'd2818401612;
        ram[249][31:0] = 32'd3198640842;
        ram[249][63:32] = 32'd2903693877;
        ram[249][95:64] = 32'd1480017882;
        ram[249][127:96] = 32'd3336666582;
        ram[250][31:0] = 32'd1375294821;
        ram[250][63:32] = 32'd2383024219;
        ram[250][95:64] = 32'd3103215630;
        ram[250][127:96] = 32'd1263697619;
        ram[251][31:0] = 32'd1342755918;
        ram[251][63:32] = 32'd1098300837;
        ram[251][95:64] = 32'd2390501042;
        ram[251][127:96] = 32'd3354638094;
        ram[252][31:0] = 32'd979321467;
        ram[252][63:32] = 32'd2054454801;
        ram[252][95:64] = 32'd894431798;
        ram[252][127:96] = 32'd3248632964;
        ram[253][31:0] = 32'd4031553092;
        ram[253][63:32] = 32'd519919884;
        ram[253][95:64] = 32'd3470978515;
        ram[253][127:96] = 32'd2062647632;
        ram[254][31:0] = 32'd595270188;
        ram[254][63:32] = 32'd3436629987;
        ram[254][95:64] = 32'd3013633939;
        ram[254][127:96] = 32'd3823758254;
        ram[255][31:0] = 32'd1993492834;
        ram[255][63:32] = 32'd707276233;
        ram[255][95:64] = 32'd401803004;
        ram[255][127:96] = 32'd1969797033;

    end
    always @(posedge clk) begin
        addr_r <= raddr;
        if(we) ram[waddr] <= din;
    end
    assign dout = ram[addr_r]; 

endmodule
